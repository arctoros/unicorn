module Unicornz_64x32 (clk, rst, arch_output_enable, arch_output_value, arch_input_enable, arch_input_value);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  output  wire [0:0] arch_output_enable;
  output  wire [7:0] arch_output_value;
  output  wire [0:0] arch_input_enable;
  input  wire [7:0] arch_input_value;

  TC_Program # (.UUID(64'd2054094413772625173 ^ UUID), .WORD_WIDTH(64'd16), .DEFAULT_FILE_NAME("Program_1C819BFC7C081515.w16.bin"), .ARG_SIG("Program_1C819BFC7C081515=%s")) Program_0 (.clk(clk), .rst(rst), .address(wire_237), .out0(wire_84), .out1(wire_225), .out2(wire_11), .out3(wire_327));
  TC_Decoder3 # (.UUID(64'd2564548179517358600 ^ UUID)) Decoder3_1 (.dis(wire_107), .sel0(wire_215), .sel1(wire_31), .sel2(wire_144), .out0(wire_87), .out1(wire_443), .out2(wire_29), .out3(wire_372), .out4(wire_474), .out5(wire_286), .out6(wire_211), .out7(wire_320));
  TC_Decoder3 # (.UUID(64'd3856915764158948127 ^ UUID)) Decoder3_2 (.dis(wire_198), .sel0(wire_215), .sel1(wire_31), .sel2(wire_144), .out0(wire_272), .out1(wire_77), .out2(wire_136), .out3(wire_329), .out4(wire_181), .out5(wire_389), .out6(wire_354), .out7(wire_171));
  TC_Decoder3 # (.UUID(64'd469263968959042607 ^ UUID)) Decoder3_3 (.dis(wire_339), .sel0(wire_215), .sel1(wire_31), .sel2(wire_144), .out0(wire_448), .out1(wire_253), .out2(wire_266), .out3(wire_167), .out4(wire_285), .out5(wire_206), .out6(wire_317), .out7(wire_278));
  TC_Decoder3 # (.UUID(64'd2355515313084503399 ^ UUID)) Decoder3_4 (.dis(wire_268), .sel0(wire_215), .sel1(wire_31), .sel2(wire_144), .out0(wire_438), .out1(wire_379), .out2(wire_202), .out3(wire_466), .out4(wire_370), .out5(wire_200), .out6(wire_456), .out7(wire_33));
  TC_Maker8 # (.UUID(64'd3412742270897961611 ^ UUID)) Maker8_5 (.in0(wire_87), .in1(wire_443), .in2(wire_29), .in3(wire_372), .in4(wire_474), .in5(wire_286), .in6(wire_211), .in7(wire_320), .out(wire_149));
  TC_Maker8 # (.UUID(64'd2545466735680713447 ^ UUID)) Maker8_6 (.in0(wire_272), .in1(wire_77), .in2(wire_136), .in3(wire_329), .in4(wire_181), .in5(wire_389), .in6(wire_354), .in7(wire_171), .out(wire_160));
  TC_Maker8 # (.UUID(64'd2498328128700172685 ^ UUID)) Maker8_7 (.in0(wire_448), .in1(wire_253), .in2(wire_266), .in3(wire_167), .in4(wire_285), .in5(wire_206), .in6(wire_317), .in7(wire_278), .out(wire_252));
  TC_Maker8 # (.UUID(64'd3307623088924666213 ^ UUID)) Maker8_8 (.in0(wire_438), .in1(wire_379), .in2(wire_202), .in3(wire_466), .in4(wire_370), .in5(wire_200), .in6(wire_456), .in7(wire_33), .out(wire_371));
  TC_Maker32 # (.UUID(64'd3223173008764962790 ^ UUID)) Maker32_9 (.in0(wire_371), .in1(wire_252), .in2(wire_160), .in3(wire_149), .out(wire_248));
  TC_Switch # (.UUID(64'd1126631217811470669 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_10 (.en(wire_449), .in(wire_21), .out(wire_47));
  TC_Switch # (.UUID(64'd383016835864160285 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_11 (.en(wire_228), .in(wire_58), .out(wire_24_0));
  TC_Switch # (.UUID(64'd3140243124393805415 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_12 (.en(wire_416), .in(wire_128), .out(wire_147));
  TC_Switch # (.UUID(64'd1581886471977480656 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_13 (.en(wire_79), .in(wire_128), .out(wire_5_0));
  TC_Switch # (.UUID(64'd2241249704231886051 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_14 (.en(wire_76), .in(wire_11[15:0]), .out(wire_58));
  TC_Switch # (.UUID(64'd4100643114395522594 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_15 (.en(wire_166), .in(wire_225[15:0]), .out(wire_21_0));
  TC_Switch # (.UUID(64'd8725165111331077 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_16 (.en(wire_146), .in(wire_11[15:0]), .out(wire_21_1));
  TC_Switch # (.UUID(64'd3499335185666676498 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_17 (.en(wire_76), .in(wire_327[15:0]), .out(wire_21_2));
  TC_And3 # (.UUID(64'd2537048141319315915 ^ UUID), .BIT_WIDTH(64'd1)) And3_18 (.in0(wire_19), .in1(wire_176), .in2(wire_159), .out(wire_175));
  TC_Program # (.UUID(64'd388994960009383908 ^ UUID), .WORD_WIDTH(64'd32), .DEFAULT_FILE_NAME("Program_565FCDAEAC6CFE4.w32.bin"), .ARG_SIG("Program_565FCDAEAC6CFE4=%s")) Program_19 (.clk(clk), .rst(rst), .address({{8{1'b0}}, wire_157 }), .out0(wire_113), .out1(), .out2(), .out3());
  TC_Not # (.UUID(64'd2992010998666944854 ^ UUID), .BIT_WIDTH(64'd1)) Not_20 (.in(wire_172), .out(wire_445));
  TC_Switch # (.UUID(64'd92717477479612822 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_21 (.en(wire_430), .in(wire_57), .out(wire_152));
  TC_Counter # (.UUID(64'd388538542796967315 ^ UUID), .BIT_WIDTH(64'd16), .count(16'd1)) Counter16_22 (.clk(clk), .rst(rst), .save(wire_172), .in(wire_125), .out(wire_387));
  TC_Counter # (.UUID(64'd3159443906265585347 ^ UUID), .BIT_WIDTH(64'd16), .count(16'd1)) Counter16_23 (.clk(clk), .rst(rst), .save(wire_60), .in(wire_125), .out(wire_36));
  TC_DelayLine # (.UUID(64'd1367561201104940128 ^ UUID), .BIT_WIDTH(64'd16)) DelayLine16_24 (.clk(clk), .rst(rst), .in(wire_15[15:0]), .out(wire_57));
  TC_Switch # (.UUID(64'd4093327232412684622 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_25 (.en(wire_172), .in(wire_36), .out(wire_97_0));
  TC_Switch # (.UUID(64'd3521663283135285715 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_26 (.en(wire_445), .in(wire_387), .out(wire_97_1));
  TC_Mux # (.UUID(64'd3040671060942591441 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_27 (.sel(wire_430), .in0(wire_97), .in1(wire_152), .out(wire_237));
  TC_DelayLine # (.UUID(64'd1970975974056862148 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_28 (.clk(clk), .rst(rst), .in(wire_2), .out(wire_430));
  TC_DelayLine # (.UUID(64'd4083747472069111906 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_29 (.clk(clk), .rst(rst), .in(wire_172), .out(wire_60));
  TC_Not # (.UUID(64'd2703499132143664233 ^ UUID), .BIT_WIDTH(64'd1)) Not_30 (.in(wire_60), .out(wire_172));
  TC_Not # (.UUID(64'd668729040907233308 ^ UUID), .BIT_WIDTH(64'd1)) Not_31 (.in(wire_144), .out(wire_431));
  TC_Not # (.UUID(64'd1492999759409908823 ^ UUID), .BIT_WIDTH(64'd1)) Not_32 (.in(wire_215), .out(wire_201));
  TC_And3 # (.UUID(64'd3485287916682882951 ^ UUID), .BIT_WIDTH(64'd1)) And3_33 (.in0(wire_431), .in1(wire_31), .in2(wire_201), .out(wire_159));
  TC_Switch # (.UUID(64'd1180978168546894742 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_34 (.en(wire_175), .in(wire_175), .out(wire_178_2));
  TC_Switch # (.UUID(64'd3723419762929890741 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_35 (.en(wire_146), .in(wire_146), .out(wire_178_1));
  TC_Switch # (.UUID(64'd2050768528734077835 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_36 (.en(wire_76), .in(wire_76), .out(wire_178_0));
  TC_Switch # (.UUID(64'd3057161046631511266 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_37 (.en(wire_294), .in(wire_294), .out(wire_146));
  TC_Decoder2 # (.UUID(64'd3508168605160458460 ^ UUID)) Decoder2_38 (.sel0(wire_222), .sel1(wire_122), .out0(), .out1(), .out2(wire_331), .out3(wire_294));
  TC_Not # (.UUID(64'd1768466669334456870 ^ UUID), .BIT_WIDTH(64'd1)) Not_39 (.in(wire_175), .out(wire_450));
  TC_Not # (.UUID(64'd3282289532960715218 ^ UUID), .BIT_WIDTH(64'd1)) Not_40 (.in(wire_250), .out(wire_198));
  TC_Not # (.UUID(64'd1327891776776277559 ^ UUID), .BIT_WIDTH(64'd1)) Not_41 (.in(wire_383), .out(wire_339));
  TC_Not # (.UUID(64'd1982359815710823425 ^ UUID), .BIT_WIDTH(64'd1)) Not_42 (.in(wire_154), .out(wire_268));
  TC_Decoder2 # (.UUID(64'd2605064451303635720 ^ UUID)) Decoder2_43 (.sel0(wire_176), .sel1(wire_19), .out0(wire_154), .out1(wire_383), .out2(wire_250), .out3(wire_179));
  TC_Add # (.UUID(64'd3313543325696297390 ^ UUID), .BIT_WIDTH(64'd16)) Add16_44 (.in0(wire_237), .in1(wire_113[15:0]), .ci(1'd0), .out(wire_125), .co());
  TC_IndexerBit # (.UUID(64'd2196806765189308211 ^ UUID), .INDEX(64'd1)) IndexerBit_45 (.in(wire_113), .out(wire_122));
  TC_IndexerBit # (.UUID(64'd737839460036088508 ^ UUID), .INDEX(64'd0)) IndexerBit_46 (.in(wire_113), .out(wire_222));
  TC_IndexerBit # (.UUID(64'd2903462054980356400 ^ UUID), .INDEX(64'd2)) IndexerBit_47 (.in(wire_113), .out(wire_76));
  TC_Splitter8 # (.UUID(64'd3910511016620535394 ^ UUID)) Splitter8_48 (.in(wire_460), .out0(wire_95), .out1(wire_83), .out2(wire_108), .out3(wire_297), .out4(wire_141), .out5(wire_22), .out6(wire_338), .out7(wire_362));
  TC_IndexerByte # (.UUID(64'd2436263972142084427 ^ UUID), .INDEX(64'd1)) IndexerByte_49 (.in({{32{1'b0}}, wire_248 }), .out(wire_460));
  TC_Switch # (.UUID(64'd607808644696146469 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_50 (.en(wire_95), .in(wire_174), .out(wire_15_5[15:0]));
  TC_Switch # (.UUID(64'd2632353714035774615 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_51 (.en(wire_83), .in(wire_243), .out(wire_15_7[15:0]));
  TC_Switch # (.UUID(64'd2222450423847071001 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_52 (.en(wire_108), .in(wire_433), .out(wire_15_9[15:0]));
  TC_Switch # (.UUID(64'd3314256307520299439 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_53 (.en(wire_297), .in(wire_88), .out(wire_15_10[15:0]));
  TC_Switch # (.UUID(64'd2595134878720988598 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_54 (.en(wire_141), .in(wire_257), .out(wire_15_12[15:0]));
  TC_Switch # (.UUID(64'd1299382207876995858 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_55 (.en(wire_22), .in(wire_455), .out(wire_15_14[15:0]));
  TC_Switch # (.UUID(64'd1287692551111612372 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_56 (.en(wire_338), .in(wire_17), .out(wire_15_16[15:0]));
  TC_Switch # (.UUID(64'd1141911395405296382 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_57 (.en(wire_362), .in({{8{1'b0}}, wire_195 }), .out(wire_15_17[15:0]));
  TC_Not # (.UUID(64'd3575339823787626444 ^ UUID), .BIT_WIDTH(64'd8)) Not8_58 (.in(wire_5[7:0]), .out(wire_195));
  TC_Rol # (.UUID(64'd2078177537373562034 ^ UUID), .BIT_WIDTH(64'd16)) Rol16_59 (.in(wire_5), .shift(wire_24[7:0]), .out(wire_17));
  TC_Shl # (.UUID(64'd4491813690601887022 ^ UUID), .BIT_WIDTH(64'd16)) Shl16_60 (.in(wire_5), .shift(wire_24[7:0]), .out(wire_257));
  TC_Shr # (.UUID(64'd4199576277751456538 ^ UUID), .BIT_WIDTH(64'd16)) Shr16_61 (.in(wire_5), .shift(wire_24[7:0]), .out(wire_88));
  TC_Xor # (.UUID(64'd1780129286836567965 ^ UUID), .BIT_WIDTH(64'd16)) Xor16_62 (.in0(wire_5), .in1(wire_24), .out(wire_433));
  TC_Or # (.UUID(64'd3629729579801707084 ^ UUID), .BIT_WIDTH(64'd16)) Or16_63 (.in0(wire_5), .in1(wire_24), .out(wire_243));
  TC_And # (.UUID(64'd3161317497787028707 ^ UUID), .BIT_WIDTH(64'd16)) And16_64 (.in0(wire_5), .in1(wire_24), .out(wire_174));
  TC_And # (.UUID(64'd381639147620396883 ^ UUID), .BIT_WIDTH(64'd8)) And8_65 (.in0(wire_304), .in1(wire_84[7:0]), .out(wire_157));
  TC_Or3 # (.UUID(64'd3488800466009071346 ^ UUID), .BIT_WIDTH(64'd1)) Or3_66 (.in0(wire_220), .in1(wire_120), .in2(wire_182), .out(wire_439));
  TC_Or # (.UUID(64'd800125638954551844 ^ UUID), .BIT_WIDTH(64'd1)) Or_67 (.in0(wire_183), .in1(wire_120), .out(wire_427));
  TC_Neg # (.UUID(64'd3923101654540497550 ^ UUID), .BIT_WIDTH(64'd16)) Neg16_68 (.in(wire_104), .out(wire_357));
  TC_Mux # (.UUID(64'd4466247896286800046 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_69 (.sel(wire_283), .in0(wire_357), .in1(wire_104), .out(wire_407));
  TC_Mux # (.UUID(64'd4573628848997923160 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_70 (.sel(wire_126), .in0({{8{1'b0}}, wire_428 }), .in1(wire_24), .out(wire_92));
  TC_Ashr # (.UUID(64'd2002805807653529301 ^ UUID), .BIT_WIDTH(64'd16)) Ashr16_71 (.in(wire_5), .shift(wire_24[7:0]), .out(wire_229));
  TC_Neg # (.UUID(64'd1410727121580829106 ^ UUID), .BIT_WIDTH(64'd16)) Neg16_72 (.in(wire_5), .out(wire_392));
  TC_Mul # (.UUID(64'd409697540344457906 ^ UUID), .BIT_WIDTH(64'd16)) DivMod16_73 (.in0(wire_5), .in1(wire_92), .out0(wire_52), .out1());
  TC_Mul # (.UUID(64'd4230356226461292418 ^ UUID), .BIT_WIDTH(64'd16)) Mul16_74 (.in0(wire_24), .in1(wire_5), .out0(wire_124), .out1());
  TC_Add # (.UUID(64'd1348307715225101930 ^ UUID), .BIT_WIDTH(64'd16)) Add16_75 (.in0(wire_407), .in1(wire_5), .ci(1'd0), .out(wire_112), .co());
  TC_Switch # (.UUID(64'd3604076901724081385 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_76 (.en(wire_0), .in(wire_392), .out(wire_15_0[15:0]));
  TC_Switch # (.UUID(64'd4522803089722429170 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_77 (.en(wire_126), .in(wire_52), .out(wire_15_2[15:0]));
  TC_Switch # (.UUID(64'd202434256468217393 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_78 (.en(wire_39), .in(wire_124), .out(wire_15_3[15:0]));
  TC_Switch # (.UUID(64'd981527730647914060 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_79 (.en(wire_439), .in(wire_112), .out(wire_15_4[15:0]));
  TC_IndexerByte # (.UUID(64'd4236276122307665751 ^ UUID), .INDEX(64'd0)) IndexerByte_80 (.in({{32{1'b0}}, wire_248 }), .out(wire_299));
  TC_Splitter8 # (.UUID(64'd4515369816812696921 ^ UUID)) Splitter8_81 (.in(wire_299), .out0(wire_182), .out1(wire_120), .out2(wire_39), .out3(wire_126), .out4(wire_0), .out5(wire_324), .out6(wire_183), .out7(wire_298));
  TC_Or # (.UUID(64'd3775589699623562439 ^ UUID), .BIT_WIDTH(64'd1)) Or_82 (.in0(wire_324), .in1(wire_183), .out(wire_220));
  TC_Or # (.UUID(64'd119900405875326486 ^ UUID), .BIT_WIDTH(64'd1)) Or_83 (.in0(wire_289), .in1(wire_114), .out(wire_138));
  TC_Add # (.UUID(64'd2771599484257026352 ^ UUID), .BIT_WIDTH(64'd16)) Add16_84 (.in0(wire_280), .in1(wire_373), .ci(1'd0), .out(wire_290), .co());
  TC_Mux # (.UUID(64'd1916750704823682311 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_85 (.sel(wire_23), .in0(wire_219), .in1(wire_47), .out(wire_282));
  TC_Switch # (.UUID(64'd110187611622282684 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_86 (.en(wire_28), .in(wire_315[15:0]), .out(wire_24_1));
  TC_Or # (.UUID(64'd1550338206798762433 ^ UUID), .BIT_WIDTH(64'd1)) Or_87 (.in0(wire_74), .in1(wire_30), .out(wire_35));
  TC_Switch # (.UUID(64'd1104805846581678264 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_88 (.en(wire_35), .in(wire_38[15:0]), .out(wire_5_1));
  TC_Or # (.UUID(64'd1973201053711173902 ^ UUID), .BIT_WIDTH(64'd1)) Or_89 (.in0(wire_30), .in1(wire_150), .out(wire_276));
  TC_And # (.UUID(64'd373051892767174731 ^ UUID), .BIT_WIDTH(64'd1)) And_90 (.in0(wire_221), .in1(wire_74), .out(wire_150));
  TC_Mux # (.UUID(64'd2189639269723513602 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_91 (.sel(wire_221), .in0(wire_336), .in1(wire_125), .out(wire_386));
  TC_Or3 # (.UUID(64'd4386189682368290849 ^ UUID), .BIT_WIDTH(64'd1)) Or3_92 (.in0(wire_30), .in1(wire_269), .in2(wire_221), .out(wire_457));
  TC_Nor # (.UUID(64'd3810192346818398090 ^ UUID), .BIT_WIDTH(64'd1)) Nor_93 (.in0(wire_457), .in1(wire_7), .out(wire_90));
  TC_Mux # (.UUID(64'd4107077995071586514 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_94 (.sel(wire_90), .in0(wire_386), .in1(wire_15[15:0]), .out(wire_177));
  TC_Switch # (.UUID(64'd1346494715147404059 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_95 (.en(wire_292), .in(wire_265), .out(wire_2_2));
  TC_Splitter8 # (.UUID(64'd3709071160935573773 ^ UUID)) Splitter8_96 (.in(wire_340), .out0(wire_41), .out1(wire_305), .out2(wire_109), .out3(wire_69), .out4(wire_300), .out5(wire_191), .out6(wire_292), .out7(wire_245));
  TC_Switch # (.UUID(64'd4272543595848591881 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_97 (.en(wire_305), .in(wire_40), .out(wire_2_7));
  TC_Switch # (.UUID(64'd2673250751246411725 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_98 (.en(wire_109), .in(wire_310), .out(wire_2_6));
  TC_Switch # (.UUID(64'd4158444071236719644 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_99 (.en(wire_69), .in(wire_472), .out(wire_2_5));
  TC_Switch # (.UUID(64'd1076960299062071464 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_100 (.en(wire_300), .in(wire_49), .out(wire_2_4));
  TC_Switch # (.UUID(64'd2871129963461955678 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_101 (.en(wire_191), .in(wire_314), .out(wire_2_3));
  TC_Switch # (.UUID(64'd1466219000736428262 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_102 (.en(wire_245), .in(wire_330), .out(wire_2_1));
  TC_LessU # (.UUID(64'd70784060852193480 ^ UUID), .BIT_WIDTH(64'd16)) LessU16_103 (.in0(wire_24), .in1(wire_5), .out(wire_330));
  TC_Or # (.UUID(64'd2633850717105506955 ^ UUID), .BIT_WIDTH(64'd1)) Or_104 (.in0(wire_330), .in1(wire_49), .out(wire_265));
  TC_Not # (.UUID(64'd2994142474806724920 ^ UUID), .BIT_WIDTH(64'd1)) Not_105 (.in(wire_49), .out(wire_314));
  TC_Equal # (.UUID(64'd4180772301230732474 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_106 (.in0(wire_5), .in1(wire_24), .out(wire_49));
  TC_LessU # (.UUID(64'd3216607671565821129 ^ UUID), .BIT_WIDTH(64'd16)) LessU16_107 (.in0(wire_5), .in1(wire_24), .out(wire_310));
  TC_Or # (.UUID(64'd1733367887190953979 ^ UUID), .BIT_WIDTH(64'd1)) Or_108 (.in0(wire_49), .in1(wire_310), .out(wire_472));
  TC_Equal # (.UUID(64'd2756161344151621510 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_109 (.in0({{8{1'b0}}, wire_214 }), .in1(wire_5), .out(wire_93));
  TC_Constant # (.UUID(64'd14059539423913175 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h0)) Constant8_110 (.out(wire_214));
  TC_Not # (.UUID(64'd2912282656104074477 ^ UUID), .BIT_WIDTH(64'd1)) Not_111 (.in(wire_93), .out(wire_40));
  TC_Switch # (.UUID(64'd338503895939097385 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_112 (.en(wire_41), .in(wire_93), .out(wire_2_8));
  TC_Switch # (.UUID(64'd2974250978505416008 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_113 (.en(wire_7), .in(wire_5), .out(wire_336));
  TC_Switch # (.UUID(64'd294942412853573551 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_114 (.en(wire_334), .in(wire_118), .out(wire_143_1));
  TC_Switch # (.UUID(64'd2530020128287448865 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_115 (.en(wire_429), .in(wire_186), .out(wire_143_0));
  TC_Not # (.UUID(64'd1944022449022311076 ^ UUID), .BIT_WIDTH(64'd1)) Not_116 (.in(wire_334), .out(wire_429));
  TC_Switch # (.UUID(64'd640117511591385720 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_117 (.en(wire_276), .in(wire_5), .out(wire_15_8[15:0]));
  TC_Clock # (.UUID(64'd473244454118914110 ^ UUID)) Clock_118 (.clk(clk), .rst(rst), .out(wire_334));
  TC_Switch # (.UUID(64'd3240978896697767469 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_119 (.en(wire_32), .in(wire_32), .out(wire_2_9));
  TC_Mux # (.UUID(64'd4327728578462997473 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_120 (.sel(wire_114), .in0(wire_282), .in1(wire_290), .out(wire_186));
  TC_Not # (.UUID(64'd2335834251709147674 ^ UUID), .BIT_WIDTH(64'd1)) Not_121 (.in(wire_258), .out(wire_449));
  TC_Switch # (.UUID(64'd1177966569030928993 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_122 (.en(wire_258), .in(wire_21), .out(wire_15_6[15:0]));
  TC_Switch # (.UUID(64'd4085565154656183842 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_123 (.en(wire_298), .in(wire_229), .out(wire_15_1[15:0]));
  TC_IndexerByte # (.UUID(64'd82359665637793120 ^ UUID), .INDEX(64'd2)) IndexerByte_124 (.in({{32{1'b0}}, wire_248 }), .out(wire_340));
  TC_Switch # (.UUID(64'd691486037870060392 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_125 (.en(wire_444), .in(wire_58), .out(wire_227));
  TC_IndexerBit # (.UUID(64'd1630189301439907508 ^ UUID), .INDEX(64'd4)) IndexerBit_126 (.in({{56{1'b0}}, wire_163 }), .out(wire_23));
  TC_IndexerBit # (.UUID(64'd2208263359456905046 ^ UUID), .INDEX(64'd5)) IndexerBit_127 (.in({{56{1'b0}}, wire_163 }), .out(wire_66));
  TC_IndexerByte # (.UUID(64'd2160584388702904456 ^ UUID), .INDEX(64'd3)) IndexerByte_128 (.in({{32{1'b0}}, wire_248 }), .out(wire_163));
  TC_Not # (.UUID(64'd904891828379418593 ^ UUID), .BIT_WIDTH(64'd1)) Not_129 (.in(wire_66), .out(wire_233));
  TC_Constant # (.UUID(64'd3538634162844758805 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hFF)) Constant8_130 (.out(wire_381));
  TC_Constant # (.UUID(64'd2648359173322761393 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hFE)) Constant8_131 (.out(wire_224));
  TC_Maker16 # (.UUID(64'd4168581648613032575 ^ UUID)) Maker16_132 (.in0(wire_381), .in1(wire_224), .out(wire_382));
  TC_Mux # (.UUID(64'd3090540701337537666 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_133 (.sel(wire_289), .in0(wire_390), .in1(wire_290), .out(wire_118));
  TC_Maker16 # (.UUID(64'd851087207377417069 ^ UUID)) Maker16_134 (.in0(wire_205), .in1(wire_420), .out(wire_373));
  TC_Constant # (.UUID(64'd381873739773538407 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hFF)) Constant8_135 (.out(wire_205));
  TC_Mux # (.UUID(64'd4592224200207251913 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_136 (.sel(wire_233), .in0(wire_73), .in1(wire_147), .out(wire_219));
  TC_Equal # (.UUID(64'd3099658865939077738 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_137 (.in0(wire_227), .in1(16'd0), .out(wire_270));
  TC_Not # (.UUID(64'd4471125710935676612 ^ UUID), .BIT_WIDTH(64'd1)) Not_138 (.in(wire_270), .out(wire_28));
  TC_IndexerBit # (.UUID(64'd460606693629125729 ^ UUID), .INDEX(64'd4)) IndexerBit_139 (.in({{56{1'b0}}, wire_153 }), .out(wire_221));
  TC_IndexerBit # (.UUID(64'd1499309531990315318 ^ UUID), .INDEX(64'd1)) IndexerBit_140 (.in({{56{1'b0}}, wire_153 }), .out(wire_269));
  TC_Or3 # (.UUID(64'd3834216222200410896 ^ UUID), .BIT_WIDTH(64'd1)) Or3_141 (.in0(wire_311), .in1(wire_325), .in2(wire_359), .out(wire_7));
  TC_IndexerBit # (.UUID(64'd345801079655292532 ^ UUID), .INDEX(64'd2)) IndexerBit_142 (.in({{56{1'b0}}, wire_153 }), .out(wire_325));
  TC_IndexerBit # (.UUID(64'd3857678701898454921 ^ UUID), .INDEX(64'd3)) IndexerBit_143 (.in({{56{1'b0}}, wire_153 }), .out(wire_311));
  TC_IndexerBit # (.UUID(64'd1094550749412879412 ^ UUID), .INDEX(64'd5)) IndexerBit_144 (.in({{56{1'b0}}, wire_153 }), .out(wire_30));
  TC_Not # (.UUID(64'd295801019876953925 ^ UUID), .BIT_WIDTH(64'd1)) Not_145 (.in(wire_179), .out(wire_107));
  TC_Equal # (.UUID(64'd3140328761418953014 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_146 (.in0(wire_118), .in1(16'd0), .out(wire_271));
  TC_Not # (.UUID(64'd4400946405007906585 ^ UUID), .BIT_WIDTH(64'd1)) Not_147 (.in(wire_440), .out(wire_74));
  TC_IndexerByte # (.UUID(64'd2633087214037843825 ^ UUID), .INDEX(64'd3)) IndexerByte_148 (.in({{32{1'b0}}, wire_248 }), .out(wire_153));
  TC_Equal # (.UUID(64'd2561182539117830921 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_149 (.in0(16'd0), .in1(wire_186), .out(wire_440));
  TC_IndexerBit # (.UUID(64'd2047893359182210890 ^ UUID), .INDEX(64'd0)) IndexerBit_150 (.in(wire_84), .out(wire_215));
  TC_IndexerBit # (.UUID(64'd3859884203355858265 ^ UUID), .INDEX(64'd1)) IndexerBit_151 (.in(wire_84), .out(wire_31));
  TC_IndexerBit # (.UUID(64'd4287739567158645737 ^ UUID), .INDEX(64'd2)) IndexerBit_152 (.in(wire_84), .out(wire_144));
  TC_IndexerBit # (.UUID(64'd777253982648504148 ^ UUID), .INDEX(64'd3)) IndexerBit_153 (.in(wire_84), .out(wire_176));
  TC_IndexerBit # (.UUID(64'd1771789865896455183 ^ UUID), .INDEX(64'd4)) IndexerBit_154 (.in(wire_84), .out(wire_19));
  TC_IndexerBit # (.UUID(64'd3105812192345802732 ^ UUID), .INDEX(64'd6)) IndexerBit_155 (.in(wire_84), .out(wire_228));
  TC_IndexerBit # (.UUID(64'd3077471030622112266 ^ UUID), .INDEX(64'd7)) IndexerBit_156 (.in(wire_84), .out(wire_79));
  TC_Not # (.UUID(64'd2159748274689718655 ^ UUID), .BIT_WIDTH(64'd1)) Not_157 (.in(wire_271), .out(wire_451));
  TC_Splitter16 # (.UUID(64'd1069070463351244943 ^ UUID)) Splitter16_158 (.in(wire_84[15:0]), .out0(), .out1(wire_332));
  TC_Switch # (.UUID(64'd3542778498052595836 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_159 (.en(wire_302), .in(wire_343[15:0]), .out(wire_15_18[15:0]));
  TC_Not # (.UUID(64'd944680686405816927 ^ UUID), .BIT_WIDTH(64'd1)) Not_160 (.in(wire_106), .out(wire_131));
  TC_Switch # (.UUID(64'd816465745217087424 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_161 (.en(wire_72), .in(wire_24), .out(wire_13));
  TC_Switch # (.UUID(64'd209623535459112064 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_162 (.en(wire_72), .in(wire_5), .out(wire_6));
  TC_And # (.UUID(64'd2522855677877010919 ^ UUID), .BIT_WIDTH(64'd1)) And_163 (.in0(wire_72), .in1(wire_437), .out(wire_302));
  TC_Equal # (.UUID(64'd2756262866884777429 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_164 (.in0(8'd0), .in1(wire_6[7:0]), .out(wire_437));
  TC_Equal # (.UUID(64'd1714264829042601315 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_165 (.in0(wire_332), .in1(wire_446), .out(wire_72));
  TC_Constant # (.UUID(64'd2907468583675662890 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_166 (.out(wire_446));
  TC_Mux # (.UUID(64'd2441497898305995710 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_167 (.sel(wire_23), .in0(wire_47), .in1(wire_73), .out(wire_390));
  TC_Switch # (.UUID(64'd3809517357945142409 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_168 (.en(wire_178), .in(wire_225[15:0]), .out(wire_128));
  TC_Not # (.UUID(64'd4003951151984714090 ^ UUID), .BIT_WIDTH(64'd1)) Not_169 (.in(wire_79), .out(wire_416));
  TC_IndexerBit # (.UUID(64'd1553590145675495351 ^ UUID), .INDEX(64'd5)) IndexerBit_170 (.in(wire_84), .out(wire_258));
  TC_Not # (.UUID(64'd3312304652180753239 ^ UUID), .BIT_WIDTH(64'd1)) Not_171 (.in(wire_228), .out(wire_444));
  TC_Constant # (.UUID(64'd2729531845625831067 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_172 (.out(wire_428));
  TC_Not # (.UUID(64'd2538698523318428916 ^ UUID), .BIT_WIDTH(64'd1)) Not_173 (.in(wire_427), .out(wire_283));
  TC_Constant # (.UUID(64'd2179489257373318160 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_174 (.out(wire_197));
  TC_Mux # (.UUID(64'd2429066787419951843 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_175 (.sel(wire_220), .in0(wire_24), .in1({{8{1'b0}}, wire_197 }), .out(wire_104));
  TC_Switch # (.UUID(64'd391371808230282023 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_176 (.en(wire_450), .in(wire_331), .out(wire_166));
  TC_Constant # (.UUID(64'd2691125905525222303 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1F)) Constant8_177 (.out(wire_304));
  TC_IndexerByte # (.UUID(64'd2112170900386343144 ^ UUID), .INDEX(64'd3)) IndexerByte_178 (.in({{32{1'b0}}, wire_248 }), .out(wire_352));
  TC_IndexerBit # (.UUID(64'd2727080739164391000 ^ UUID), .INDEX(64'd6)) IndexerBit_179 (.in({{56{1'b0}}, wire_352 }), .out(wire_1));
  TC_Switch # (.UUID(64'd2160087561000370162 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_180 (.en(wire_1), .in(wire_1), .out(wire_2_0));
  TC_Switch # (.UUID(64'd592302940647155691 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_181 (.en(wire_242), .in({{15{1'b0}}, wire_34 }), .out(wire_15_11[15:0]));
  TC_Or # (.UUID(64'd3278179513885088927 ^ UUID), .BIT_WIDTH(64'd1)) Or_182 (.in0(wire_242), .in1(wire_100), .out(wire_296));
  TC_Equal # (.UUID(64'd4033274235037801114 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_183 (.in0(wire_471), .in1(wire_99), .out(wire_242));
  TC_Not # (.UUID(64'd1697593568395826930 ^ UUID), .BIT_WIDTH(64'd1)) Not_184 (.in(wire_100), .out(wire_85));
  TC_Splitter16 # (.UUID(64'd962308306064647197 ^ UUID)) Splitter16_185 (.in(wire_84[15:0]), .out0(), .out1(wire_471));
  TC_Constant # (.UUID(64'd3037869375563223000 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h2)) Constant8_186 (.out(wire_99));
  TC_DelayLine # (.UUID(64'd4275385609773382257 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_187 (.clk(clk), .rst(rst), .in(wire_409), .out(wire_100));
  TC_Switch # (.UUID(64'd1286392688347840013 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_188 (.en(wire_85), .in(wire_296), .out(wire_409));
  TC_Splitter16 # (.UUID(64'd815166994044352782 ^ UUID)) Splitter16_189 (.in(wire_84[15:0]), .out0(), .out1(wire_261));
  TC_IndexerByte # (.UUID(64'd4056757385308142069 ^ UUID), .INDEX(64'd1)) IndexerByte_190 (.in(wire_293), .out(wire_350));
  TC_IndexerByte # (.UUID(64'd4445007758314830950 ^ UUID), .INDEX(64'd0)) IndexerByte_191 (.in(wire_293), .out(wire_421));
  TC_Maker16 # (.UUID(64'd1879612468053834457 ^ UUID)) Maker16_192 (.in0(wire_421), .in1(wire_350), .out(wire_137));
  TC_Switch # (.UUID(64'd220823607166135876 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_193 (.en(wire_365), .in(wire_137), .out(wire_15_15[15:0]));
  TC_Equal # (.UUID(64'd3724760983101447498 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_194 (.in0(wire_261), .in1(wire_369), .out(wire_365));
  TC_Constant # (.UUID(64'd1337227511337026411 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h3)) Constant8_195 (.out(wire_369));
  TC_Timing # (.UUID(64'd2799049267103079424 ^ UUID)) Timing_196 (.en(wire_365), .out(wire_293));
  TC_DotMatrixDisplay # (.UUID(64'd3664136990544334169 ^ UUID)) DotMatrixDisplay_197 (.clk(clk), .rst(rst), .en_y(wire_117[0:0]), .en_x(wire_111[0:0]), .color_info(wire_117), .pixel_info(wire_111));
  TC_DotMatrixDisplay # (.UUID(64'd4523285523904489011 ^ UUID)) DotMatrixDisplay_198 (.clk(clk), .rst(rst), .en_y(wire_27[0:0]), .en_x(wire_111[0:0]), .color_info(wire_27), .pixel_info(wire_111));
  TC_DotMatrixDisplay # (.UUID(64'd2454247312537554172 ^ UUID)) DotMatrixDisplay_199 (.clk(clk), .rst(rst), .en_y(wire_45[0:0]), .en_x(wire_111[0:0]), .color_info(wire_45), .pixel_info(wire_111));
  TC_DotMatrixDisplay # (.UUID(64'd1716960261624563378 ^ UUID)) DotMatrixDisplay_200 (.clk(clk), .rst(rst), .en_y(wire_98[0:0]), .en_x(wire_111[0:0]), .color_info(wire_98), .pixel_info(wire_111));
  TC_DotMatrixDisplay # (.UUID(64'd477724403087111064 ^ UUID)) DotMatrixDisplay_201 (.clk(clk), .rst(rst), .en_y(wire_50[0:0]), .en_x(wire_111[0:0]), .color_info(wire_50), .pixel_info(wire_111));
  TC_DotMatrixDisplay # (.UUID(64'd233502698066449431 ^ UUID)) DotMatrixDisplay_202 (.clk(clk), .rst(rst), .en_y(wire_9[0:0]), .en_x(wire_111[0:0]), .color_info(wire_9), .pixel_info(wire_111));
  TC_DotMatrixDisplay # (.UUID(64'd2643939785681194081 ^ UUID)) DotMatrixDisplay_203 (.clk(clk), .rst(rst), .en_y(wire_68[0:0]), .en_x(wire_111[0:0]), .color_info(wire_68), .pixel_info(wire_111));
  TC_DotMatrixDisplay # (.UUID(64'd2456097156852606244 ^ UUID)) DotMatrixDisplay_204 (.clk(clk), .rst(rst), .en_y(wire_133[0:0]), .en_x(wire_111[0:0]), .color_info(wire_133), .pixel_info(wire_111));
  TC_DotMatrixDisplay # (.UUID(64'd1295657997286150516 ^ UUID)) DotMatrixDisplay_205 (.clk(clk), .rst(rst), .en_y(wire_231[0:0]), .en_x(wire_111[0:0]), .color_info(wire_231), .pixel_info(wire_111));
  TC_DotMatrixDisplay # (.UUID(64'd769058939343858260 ^ UUID)) DotMatrixDisplay_206 (.clk(clk), .rst(rst), .en_y(wire_135[0:0]), .en_x(wire_111[0:0]), .color_info(wire_135), .pixel_info(wire_111));
  TC_DotMatrixDisplay # (.UUID(64'd2258332813225485225 ^ UUID)) DotMatrixDisplay_207 (.clk(clk), .rst(rst), .en_y(wire_62[0:0]), .en_x(wire_111[0:0]), .color_info(wire_62), .pixel_info(wire_111));
  TC_DotMatrixDisplay # (.UUID(64'd1094247889656016871 ^ UUID)) DotMatrixDisplay_208 (.clk(clk), .rst(rst), .en_y(wire_117[0:0]), .en_x(wire_82[0:0]), .color_info(wire_117), .pixel_info(wire_82));
  TC_DotMatrixDisplay # (.UUID(64'd2906317122771197315 ^ UUID)) DotMatrixDisplay_209 (.clk(clk), .rst(rst), .en_y(wire_27[0:0]), .en_x(wire_82[0:0]), .color_info(wire_27), .pixel_info(wire_82));
  TC_DotMatrixDisplay # (.UUID(64'd2710556982130869271 ^ UUID)) DotMatrixDisplay_210 (.clk(clk), .rst(rst), .en_y(wire_45[0:0]), .en_x(wire_82[0:0]), .color_info(wire_45), .pixel_info(wire_82));
  TC_DotMatrixDisplay # (.UUID(64'd3820587598745411362 ^ UUID)) DotMatrixDisplay_211 (.clk(clk), .rst(rst), .en_y(wire_98[0:0]), .en_x(wire_82[0:0]), .color_info(wire_98), .pixel_info(wire_82));
  TC_DotMatrixDisplay # (.UUID(64'd636375990872542647 ^ UUID)) DotMatrixDisplay_212 (.clk(clk), .rst(rst), .en_y(wire_50[0:0]), .en_x(wire_82[0:0]), .color_info(wire_50), .pixel_info(wire_82));
  TC_DotMatrixDisplay # (.UUID(64'd3918293502762045952 ^ UUID)) DotMatrixDisplay_213 (.clk(clk), .rst(rst), .en_y(wire_9[0:0]), .en_x(wire_82[0:0]), .color_info(wire_9), .pixel_info(wire_82));
  TC_DotMatrixDisplay # (.UUID(64'd3954665317158973579 ^ UUID)) DotMatrixDisplay_214 (.clk(clk), .rst(rst), .en_y(wire_68[0:0]), .en_x(wire_82[0:0]), .color_info(wire_68), .pixel_info(wire_82));
  TC_DotMatrixDisplay # (.UUID(64'd4443983821981529472 ^ UUID)) DotMatrixDisplay_215 (.clk(clk), .rst(rst), .en_y(wire_133[0:0]), .en_x(wire_82[0:0]), .color_info(wire_133), .pixel_info(wire_82));
  TC_DotMatrixDisplay # (.UUID(64'd2971913797960446620 ^ UUID)) DotMatrixDisplay_216 (.clk(clk), .rst(rst), .en_y(wire_231[0:0]), .en_x(wire_82[0:0]), .color_info(wire_231), .pixel_info(wire_82));
  TC_DotMatrixDisplay # (.UUID(64'd984824982458035893 ^ UUID)) DotMatrixDisplay_217 (.clk(clk), .rst(rst), .en_y(wire_135[0:0]), .en_x(wire_82[0:0]), .color_info(wire_135), .pixel_info(wire_82));
  TC_DotMatrixDisplay # (.UUID(64'd370313129409463494 ^ UUID)) DotMatrixDisplay_218 (.clk(clk), .rst(rst), .en_y(wire_62[0:0]), .en_x(wire_82[0:0]), .color_info(wire_62), .pixel_info(wire_82));
  TC_DotMatrixDisplay # (.UUID(64'd1659341693991075024 ^ UUID)) DotMatrixDisplay_219 (.clk(clk), .rst(rst), .en_y(wire_117[0:0]), .en_x(wire_26[0:0]), .color_info(wire_117), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd4090442229255502662 ^ UUID)) DotMatrixDisplay_220 (.clk(clk), .rst(rst), .en_y(wire_27[0:0]), .en_x(wire_26[0:0]), .color_info(wire_27), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd2120522814468093527 ^ UUID)) DotMatrixDisplay_221 (.clk(clk), .rst(rst), .en_y(wire_45[0:0]), .en_x(wire_26[0:0]), .color_info(wire_45), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd2275199029062329834 ^ UUID)) DotMatrixDisplay_222 (.clk(clk), .rst(rst), .en_y(wire_98[0:0]), .en_x(wire_26[0:0]), .color_info(wire_98), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd1393728114345846423 ^ UUID)) DotMatrixDisplay_223 (.clk(clk), .rst(rst), .en_y(wire_50[0:0]), .en_x(wire_26[0:0]), .color_info(wire_50), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd4545002377462046516 ^ UUID)) DotMatrixDisplay_224 (.clk(clk), .rst(rst), .en_y(wire_9[0:0]), .en_x(wire_26[0:0]), .color_info(wire_9), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd2517565327759169021 ^ UUID)) DotMatrixDisplay_225 (.clk(clk), .rst(rst), .en_y(wire_68[0:0]), .en_x(wire_26[0:0]), .color_info(wire_68), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd2656861857212416788 ^ UUID)) DotMatrixDisplay_226 (.clk(clk), .rst(rst), .en_y(wire_133[0:0]), .en_x(wire_26[0:0]), .color_info(wire_133), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd276436997605160609 ^ UUID)) DotMatrixDisplay_227 (.clk(clk), .rst(rst), .en_y(wire_231[0:0]), .en_x(wire_26[0:0]), .color_info(wire_231), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd259750575459531229 ^ UUID)) DotMatrixDisplay_228 (.clk(clk), .rst(rst), .en_y(wire_135[0:0]), .en_x(wire_26[0:0]), .color_info(wire_135), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd3675714028900344906 ^ UUID)) DotMatrixDisplay_229 (.clk(clk), .rst(rst), .en_y(wire_62[0:0]), .en_x(wire_26[0:0]), .color_info(wire_62), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd221996997629957745 ^ UUID)) DotMatrixDisplay_230 (.clk(clk), .rst(rst), .en_y(wire_117[0:0]), .en_x(wire_139[0:0]), .color_info(wire_117), .pixel_info(wire_139));
  TC_DotMatrixDisplay # (.UUID(64'd2106603050357944433 ^ UUID)) DotMatrixDisplay_231 (.clk(clk), .rst(rst), .en_y(wire_98[0:0]), .en_x(wire_139[0:0]), .color_info(wire_98), .pixel_info(wire_139));
  TC_DotMatrixDisplay # (.UUID(64'd253488447841708180 ^ UUID)) DotMatrixDisplay_232 (.clk(clk), .rst(rst), .en_y(wire_50[0:0]), .en_x(wire_139[0:0]), .color_info(wire_50), .pixel_info(wire_139));
  TC_DotMatrixDisplay # (.UUID(64'd612463031464991440 ^ UUID)) DotMatrixDisplay_233 (.clk(clk), .rst(rst), .en_y(wire_9[0:0]), .en_x(wire_139[0:0]), .color_info(wire_9), .pixel_info(wire_139));
  TC_DotMatrixDisplay # (.UUID(64'd2928242032974181734 ^ UUID)) DotMatrixDisplay_234 (.clk(clk), .rst(rst), .en_y(wire_68[0:0]), .en_x(wire_139[0:0]), .color_info(wire_68), .pixel_info(wire_139));
  TC_DotMatrixDisplay # (.UUID(64'd3112334513645503701 ^ UUID)) DotMatrixDisplay_235 (.clk(clk), .rst(rst), .en_y(wire_133[0:0]), .en_x(wire_139[0:0]), .color_info(wire_133), .pixel_info(wire_139));
  TC_DotMatrixDisplay # (.UUID(64'd2438205929049834623 ^ UUID)) DotMatrixDisplay_236 (.clk(clk), .rst(rst), .en_y(wire_231[0:0]), .en_x(wire_139[0:0]), .color_info(wire_231), .pixel_info(wire_139));
  TC_DotMatrixDisplay # (.UUID(64'd2583268778611470830 ^ UUID)) DotMatrixDisplay_237 (.clk(clk), .rst(rst), .en_y(wire_135[0:0]), .en_x(wire_139[0:0]), .color_info(wire_135), .pixel_info(wire_139));
  TC_DotMatrixDisplay # (.UUID(64'd1417567905964410602 ^ UUID)) DotMatrixDisplay_238 (.clk(clk), .rst(rst), .en_y(wire_62[0:0]), .en_x(wire_139[0:0]), .color_info(wire_62), .pixel_info(wire_139));
  TC_Or # (.UUID(64'd4552406311139818817 ^ UUID), .BIT_WIDTH(64'd32)) Or32_239 (.in0({{31{1'b0}}, wire_185 }), .in1(wire_3), .out(wire_117));
  TC_Or # (.UUID(64'd4379624752864373096 ^ UUID), .BIT_WIDTH(64'd32)) Or32_240 (.in0({{31{1'b0}}, wire_366 }), .in1(wire_3), .out(wire_27));
  TC_Or # (.UUID(64'd4205159359974210151 ^ UUID), .BIT_WIDTH(64'd32)) Or32_241 (.in0({{31{1'b0}}, wire_301 }), .in1(wire_3), .out(wire_98));
  TC_Or # (.UUID(64'd3475250448327390751 ^ UUID), .BIT_WIDTH(64'd32)) Or32_242 (.in0({{31{1'b0}}, wire_169 }), .in1(wire_3), .out(wire_50));
  TC_Or # (.UUID(64'd3433362640040173500 ^ UUID), .BIT_WIDTH(64'd32)) Or32_243 (.in0({{31{1'b0}}, wire_232 }), .in1(wire_3), .out(wire_9));
  TC_Or # (.UUID(64'd221937994222578023 ^ UUID), .BIT_WIDTH(64'd32)) Or32_244 (.in0({{31{1'b0}}, wire_378 }), .in1(wire_3), .out(wire_68));
  TC_Or # (.UUID(64'd1128671621782155494 ^ UUID), .BIT_WIDTH(64'd32)) Or32_245 (.in0({{31{1'b0}}, wire_148 }), .in1(wire_3), .out(wire_133));
  TC_Or # (.UUID(64'd3489283905828808476 ^ UUID), .BIT_WIDTH(64'd32)) Or32_246 (.in0({{31{1'b0}}, wire_418 }), .in1(wire_3), .out(wire_231));
  TC_Or # (.UUID(64'd4549501439555191842 ^ UUID), .BIT_WIDTH(64'd32)) Or32_247 (.in0({{31{1'b0}}, wire_61 }), .in1(wire_3), .out(wire_135));
  TC_Or # (.UUID(64'd515760107847623846 ^ UUID), .BIT_WIDTH(64'd32)) Or32_248 (.in0({{31{1'b0}}, wire_247 }), .in1(wire_3), .out(wire_62));
  TC_Decoder3 # (.UUID(64'd2355883731160852788 ^ UUID)) Decoder3_249 (.dis(wire_121), .sel0(wire_10), .sel1(wire_86), .sel2(wire_396), .out0(wire_185), .out1(wire_366), .out2(wire_328), .out3(wire_301), .out4(wire_169), .out5(wire_232), .out6(wire_378), .out7(wire_148));
  TC_Decoder2 # (.UUID(64'd43300923688619049 ^ UUID)) Decoder2_250 (.sel0(wire_10), .sel1(wire_86), .out0(wire_213), .out1(wire_184), .out2(wire_275), .out3());
  TC_Switch # (.UUID(64'd4034663872841809180 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_251 (.en(wire_121), .in(wire_213), .out(wire_418));
  TC_Switch # (.UUID(64'd2817107100876533977 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_252 (.en(wire_121), .in(wire_184), .out(wire_61));
  TC_Or # (.UUID(64'd3774487218439831887 ^ UUID), .BIT_WIDTH(64'd64)) Or64_253 (.in0(wire_187), .in1({{63{1'b0}}, wire_67 }), .out(wire_318));
  TC_Or # (.UUID(64'd4321088425401214646 ^ UUID), .BIT_WIDTH(64'd64)) Or64_254 (.in0(wire_187), .in1({{63{1'b0}}, wire_188 }), .out(wire_333));
  TC_Or # (.UUID(64'd805663505735110387 ^ UUID), .BIT_WIDTH(64'd64)) Or64_255 (.in0(wire_187), .in1({{63{1'b0}}, wire_435 }), .out(wire_142));
  TC_Maker8 # (.UUID(64'd1899838318998446938 ^ UUID)) Maker8_256 (.in0(wire_75), .in1(wire_434), .in2(wire_432), .in3(wire_180), .in4(wire_397), .in5(wire_308), .in6(wire_452), .in7(wire_459), .out(wire_259));
  TC_Maker8 # (.UUID(64'd984839894031669175 ^ UUID)) Maker8_257 (.in0(wire_470), .in1(wire_349), .in2(wire_341), .in3(wire_351), .in4(wire_347), .in5(wire_194), .in6(wire_263), .in7(wire_463), .out(wire_8));
  TC_Maker8 # (.UUID(64'd3860204027489987942 ^ UUID)) Maker8_258 (.in0(wire_116), .in1(wire_238), .in2(wire_453), .in3(wire_426), .in4(wire_287), .in5(wire_469), .in6(wire_355), .in7(wire_279), .out(wire_65));
  TC_Maker8 # (.UUID(64'd432487347562912252 ^ UUID)) Maker8_259 (.in0(wire_422), .in1(wire_274), .in2(wire_241), .in3(wire_312), .in4(wire_244), .in5(wire_164), .in6(wire_461), .in7(wire_393), .out(wire_403));
  TC_Maker8 # (.UUID(64'd3736712824354188155 ^ UUID)) Maker8_260 (.in0(wire_204), .in1(wire_316), .in2(wire_313), .in3(wire_303), .in4(wire_103), .in5(wire_476), .in6(wire_81), .in7(wire_467), .out(wire_262));
  TC_Decoder3 # (.UUID(64'd884438583600364956 ^ UUID)) Decoder3_261 (.dis(wire_80), .sel0(wire_20), .sel1(wire_16), .sel2(wire_43), .out0(wire_75), .out1(wire_434), .out2(wire_432), .out3(wire_180), .out4(wire_397), .out5(wire_308), .out6(wire_452), .out7(wire_459));
  TC_Not # (.UUID(64'd1756422684115560108 ^ UUID), .BIT_WIDTH(64'd1)) Not_262 (.in(wire_78), .out(wire_123));
  TC_And # (.UUID(64'd1263154755327333848 ^ UUID), .BIT_WIDTH(64'd1)) And_263 (.in0(wire_398), .in1(wire_475), .out(wire_260));
  TC_And3 # (.UUID(64'd2004083645781838127 ^ UUID), .BIT_WIDTH(64'd1)) And3_264 (.in0(wire_110), .in1(wire_462), .in2(wire_260), .out(wire_78));
  TC_And3 # (.UUID(64'd1884602402787279659 ^ UUID), .BIT_WIDTH(64'd1)) And3_265 (.in0(wire_346), .in1(wire_56), .in2(wire_14), .out(wire_307));
  TC_Not # (.UUID(64'd4393826969183798925 ^ UUID), .BIT_WIDTH(64'd1)) Not_266 (.in(wire_56), .out(wire_462));
  TC_And3 # (.UUID(64'd2929028691481501737 ^ UUID), .BIT_WIDTH(64'd1)) And3_267 (.in0(wire_110), .in1(wire_170), .in2(wire_42), .out(wire_363));
  TC_And # (.UUID(64'd3980703843308468025 ^ UUID), .BIT_WIDTH(64'd1)) And_268 (.in0(wire_145), .in1(wire_216), .out(wire_42));
  TC_And3 # (.UUID(64'd3008184888437837797 ^ UUID), .BIT_WIDTH(64'd1)) And3_269 (.in0(wire_442), .in1(wire_395), .in2(wire_218), .out(wire_267));
  TC_And # (.UUID(64'd854056611492606295 ^ UUID), .BIT_WIDTH(64'd1)) And_270 (.in0(wire_145), .in1(wire_410), .out(wire_218));
  TC_And3 # (.UUID(64'd932847285064479538 ^ UUID), .BIT_WIDTH(64'd1)) And3_271 (.in0(wire_110), .in1(wire_56), .in2(wire_207), .out(wire_134));
  TC_And # (.UUID(64'd723925587366255632 ^ UUID), .BIT_WIDTH(64'd1)) And_272 (.in0(wire_361), .in1(wire_364), .out(wire_207));
  TC_And # (.UUID(64'd3997202033913493589 ^ UUID), .BIT_WIDTH(64'd1)) And_273 (.in0(wire_419), .in1(wire_406), .out(wire_14));
  TC_Not # (.UUID(64'd3837755846434102303 ^ UUID), .BIT_WIDTH(64'd1)) Not_274 (.in(wire_91), .out(wire_216));
  TC_Not # (.UUID(64'd3728171245612547644 ^ UUID), .BIT_WIDTH(64'd1)) Not_275 (.in(wire_56), .out(wire_170));
  TC_Not # (.UUID(64'd2410308471969065618 ^ UUID), .BIT_WIDTH(64'd1)) Not_276 (.in(wire_110), .out(wire_442));
  TC_Not # (.UUID(64'd820998404102950992 ^ UUID), .BIT_WIDTH(64'd1)) Not_277 (.in(wire_91), .out(wire_410));
  TC_Not # (.UUID(64'd2021565867020626441 ^ UUID), .BIT_WIDTH(64'd1)) Not_278 (.in(wire_56), .out(wire_395));
  TC_Not # (.UUID(64'd2180051592468327154 ^ UUID), .BIT_WIDTH(64'd1)) Not_279 (.in(wire_91), .out(wire_364));
  TC_Not # (.UUID(64'd1820017548761317419 ^ UUID), .BIT_WIDTH(64'd1)) Not_280 (.in(wire_145), .out(wire_361));
  TC_Not # (.UUID(64'd2145258914016335304 ^ UUID), .BIT_WIDTH(64'd1)) Not_281 (.in(wire_110), .out(wire_346));
  TC_Not # (.UUID(64'd1580884975280642426 ^ UUID), .BIT_WIDTH(64'd1)) Not_282 (.in(wire_91), .out(wire_406));
  TC_Not # (.UUID(64'd995815798857176822 ^ UUID), .BIT_WIDTH(64'd1)) Not_283 (.in(wire_145), .out(wire_419));
  TC_Not # (.UUID(64'd1957814361250160086 ^ UUID), .BIT_WIDTH(64'd1)) Not_284 (.in(wire_91), .out(wire_475));
  TC_Not # (.UUID(64'd2899922533480021322 ^ UUID), .BIT_WIDTH(64'd1)) Not_285 (.in(wire_145), .out(wire_398));
  TC_Not # (.UUID(64'd4357804555026814051 ^ UUID), .BIT_WIDTH(64'd1)) Not_286 (.in(wire_363), .out(wire_80));
  TC_Not # (.UUID(64'd925031083123060575 ^ UUID), .BIT_WIDTH(64'd1)) Not_287 (.in(wire_267), .out(wire_127));
  TC_Not # (.UUID(64'd2594386124497233616 ^ UUID), .BIT_WIDTH(64'd1)) Not_288 (.in(wire_134), .out(wire_239));
  TC_Not # (.UUID(64'd1981766396418540652 ^ UUID), .BIT_WIDTH(64'd1)) Not_289 (.in(wire_307), .out(wire_391));
  TC_Decoder3 # (.UUID(64'd2347530673898705732 ^ UUID)) Decoder3_290 (.dis(wire_127), .sel0(wire_20), .sel1(wire_16), .sel2(wire_43), .out0(wire_470), .out1(wire_349), .out2(wire_341), .out3(wire_351), .out4(wire_347), .out5(wire_194), .out6(wire_263), .out7(wire_463));
  TC_Decoder3 # (.UUID(64'd2919245333301046076 ^ UUID)) Decoder3_291 (.dis(wire_239), .sel0(wire_20), .sel1(wire_16), .sel2(wire_43), .out0(wire_116), .out1(wire_238), .out2(wire_453), .out3(wire_426), .out4(wire_287), .out5(wire_469), .out6(wire_355), .out7(wire_279));
  TC_Decoder3 # (.UUID(64'd2250913747292488162 ^ UUID)) Decoder3_292 (.dis(wire_391), .sel0(wire_20), .sel1(wire_16), .sel2(wire_43), .out0(wire_422), .out1(wire_274), .out2(wire_241), .out3(wire_312), .out4(wire_244), .out5(wire_164), .out6(wire_461), .out7(wire_393));
  TC_Decoder3 # (.UUID(64'd205315477120840980 ^ UUID)) Decoder3_293 (.dis(wire_123), .sel0(wire_20), .sel1(wire_16), .sel2(wire_43), .out0(wire_204), .out1(wire_316), .out2(wire_313), .out3(wire_303), .out4(wire_103), .out5(wire_476), .out6(wire_81), .out7(wire_467));
  TC_Maker8 # (.UUID(64'd295352228004415385 ^ UUID)) Maker8_294 (.in0(wire_212), .in1(wire_119), .in2(wire_377), .in3(wire_394), .in4(wire_18), .in5(wire_284), .in6(wire_417), .in7(wire_246), .out(wire_155));
  TC_Not # (.UUID(64'd2569473202873079078 ^ UUID), .BIT_WIDTH(64'd1)) Not_295 (.in(wire_145), .out(wire_236));
  TC_Not # (.UUID(64'd549515294479480322 ^ UUID), .BIT_WIDTH(64'd1)) Not_296 (.in(wire_91), .out(wire_281));
  TC_Decoder3 # (.UUID(64'd2217537975887549640 ^ UUID)) Decoder3_297 (.dis(wire_376), .sel0(wire_20), .sel1(wire_16), .sel2(wire_43), .out0(wire_212), .out1(wire_119), .out2(wire_377), .out3(wire_394), .out4(wire_18), .out5(wire_284), .out6(wire_417), .out7(wire_246));
  TC_And3 # (.UUID(64'd3464733780494301715 ^ UUID), .BIT_WIDTH(64'd1)) And3_298 (.in0(wire_189), .in1(wire_96), .in2(wire_162), .out(wire_89));
  TC_And3 # (.UUID(64'd3673302305383611256 ^ UUID), .BIT_WIDTH(64'd1)) And3_299 (.in0(wire_399), .in1(wire_236), .in2(wire_281), .out(wire_162));
  TC_Maker64 # (.UUID(64'd2796473728191387387 ^ UUID)) Maker64_300 (.in0(8'd0), .in1(wire_155), .in2(wire_262), .in3(wire_403), .in4(wire_65), .in5(wire_8), .in6(wire_259), .in7(8'd0), .out(wire_187));
  TC_Constant # (.UUID(64'd476599345246060721 ^ UUID), .BIT_WIDTH(64'd64), .value(64'h100000000000000)) Constant64_301 (.out(wire_140));
  TC_Decoder2 # (.UUID(64'd719562623271464916 ^ UUID)) Decoder2_302 (.sel0(wire_400), .sel1(wire_408), .out0(wire_67), .out1(wire_188), .out2(wire_380), .out3(wire_435));
  TC_Or # (.UUID(64'd3933533332118879027 ^ UUID), .BIT_WIDTH(64'd64)) Or64_303 (.in0(wire_187), .in1({{63{1'b0}}, wire_380 }), .out(wire_414));
  TC_Or # (.UUID(64'd3885849532696548888 ^ UUID), .BIT_WIDTH(64'd64)) Or64_304 (.in0(wire_414), .in1(wire_140), .out(wire_26));
  TC_Or # (.UUID(64'd2771931884579429156 ^ UUID), .BIT_WIDTH(64'd64)) Or64_305 (.in0(wire_142), .in1(wire_140), .out(wire_139));
  TC_Or # (.UUID(64'd1895393282243127434 ^ UUID), .BIT_WIDTH(64'd64)) Or64_306 (.in0(wire_333), .in1(wire_140), .out(wire_82));
  TC_Or # (.UUID(64'd2126784000832456339 ^ UUID), .BIT_WIDTH(64'd64)) Or64_307 (.in0(wire_318), .in1(wire_140), .out(wire_111));
  TC_Not # (.UUID(64'd1813774519689494074 ^ UUID), .BIT_WIDTH(64'd1)) Not_308 (.in(wire_56), .out(wire_399));
  TC_IndexerBit # (.UUID(64'd4483867977540107476 ^ UUID), .INDEX(64'd0)) IndexerBit_309 (.in({{56{1'b0}}, wire_249 }), .out(wire_20));
  TC_IndexerBit # (.UUID(64'd1265819950009573605 ^ UUID), .INDEX(64'd1)) IndexerBit_310 (.in({{56{1'b0}}, wire_249 }), .out(wire_16));
  TC_IndexerBit # (.UUID(64'd3730218088294752693 ^ UUID), .INDEX(64'd2)) IndexerBit_311 (.in({{56{1'b0}}, wire_249 }), .out(wire_43));
  TC_IndexerBit # (.UUID(64'd3379558781261549428 ^ UUID), .INDEX(64'd3)) IndexerBit_312 (.in({{56{1'b0}}, wire_249 }), .out(wire_110));
  TC_IndexerBit # (.UUID(64'd2333701187965543463 ^ UUID), .INDEX(64'd4)) IndexerBit_313 (.in({{56{1'b0}}, wire_249 }), .out(wire_56));
  TC_IndexerBit # (.UUID(64'd681828137790676581 ^ UUID), .INDEX(64'd5)) IndexerBit_314 (.in({{56{1'b0}}, wire_249 }), .out(wire_145));
  TC_Maker8 # (.UUID(64'd965647765177340792 ^ UUID)) Maker8_315 (.in0(wire_12), .in1(wire_94), .in2(wire_59), .in3(wire_54), .in4(wire_12), .in5(wire_94), .in6(wire_59), .in7(wire_54), .out(wire_424));
  TC_Maker8 # (.UUID(64'd1370718817211265218 ^ UUID)) Maker8_316 (.in0(wire_240), .in1(wire_64), .in2(wire_59), .in3(wire_54), .in4(wire_240), .in5(wire_64), .in6(wire_59), .in7(wire_54), .out(wire_436));
  TC_Maker8 # (.UUID(64'd4524398156080664253 ^ UUID)) Maker8_317 (.in0(wire_368), .in1(wire_51), .in2(wire_59), .in3(wire_54), .in4(wire_368), .in5(wire_51), .in6(wire_59), .in7(wire_54), .out(wire_356));
  TC_Switch # (.UUID(64'd36275008520620059 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_318 (.en(wire_367[0:0]), .in(wire_424), .out(wire_323));
  TC_Switch # (.UUID(64'd2752121200656840932 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_319 (.en(wire_412[0:0]), .in(wire_436), .out(wire_254));
  TC_Switch # (.UUID(64'd2522875977552864454 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_320 (.en(wire_374[0:0]), .in(wire_356), .out(wire_345));
  TC_Maker32 # (.UUID(64'd4438245501521141190 ^ UUID)) Maker32_321 (.in0(8'd0), .in1(wire_345), .in2(wire_254), .in3(wire_323), .out(wire_3));
  TC_IndexerBit # (.UUID(64'd2773381416993893124 ^ UUID), .INDEX(64'd0)) IndexerBit_322 (.in({{56{1'b0}}, wire_168 }), .out(wire_12));
  TC_IndexerBit # (.UUID(64'd580753202887096457 ^ UUID), .INDEX(64'd1)) IndexerBit_323 (.in({{56{1'b0}}, wire_168 }), .out(wire_94));
  TC_IndexerBit # (.UUID(64'd1607506216411020602 ^ UUID), .INDEX(64'd2)) IndexerBit_324 (.in({{56{1'b0}}, wire_168 }), .out(wire_240));
  TC_IndexerBit # (.UUID(64'd339327870727800916 ^ UUID), .INDEX(64'd3)) IndexerBit_325 (.in({{56{1'b0}}, wire_168 }), .out(wire_64));
  TC_IndexerBit # (.UUID(64'd538049426750639330 ^ UUID), .INDEX(64'd4)) IndexerBit_326 (.in({{56{1'b0}}, wire_168 }), .out(wire_368));
  TC_IndexerBit # (.UUID(64'd3988667738118775649 ^ UUID), .INDEX(64'd5)) IndexerBit_327 (.in({{56{1'b0}}, wire_168 }), .out(wire_51));
  TC_Splitter32 # (.UUID(64'd2215188549689077647 ^ UUID)) Splitter32_328 (.in(wire_129), .out0(), .out1(wire_374), .out2(wire_412), .out3(wire_367));
  TC_Maker64 # (.UUID(64'd3058259462461040721 ^ UUID)) Maker64_329 (.in0({{7{1'b0}}, wire_12 }), .in1({{7{1'b0}}, wire_94 }), .in2({{7{1'b0}}, wire_240 }), .in3({{7{1'b0}}, wire_64 }), .in4({{7{1'b0}}, wire_368 }), .in5({{7{1'b0}}, wire_51 }), .in6(8'd0), .in7(8'd0), .out(wire_130));
  TC_Maker32 # (.UUID(64'd4302620568193657741 ^ UUID)) Maker32_330 (.in0(8'd0), .in1(wire_192), .in2(wire_226), .in3(wire_342), .out(wire_129));
  TC_Or # (.UUID(64'd803353250254897789 ^ UUID), .BIT_WIDTH(64'd8)) Or8_331 (.in0(wire_404), .in1(wire_425), .out(wire_192));
  TC_IndexerByte # (.UUID(64'd2441854781662376807 ^ UUID), .INDEX(64'd4)) IndexerByte_332 (.in(wire_130), .out(wire_404));
  TC_IndexerByte # (.UUID(64'd862882653762759736 ^ UUID), .INDEX(64'd5)) IndexerByte_333 (.in(wire_130), .out(wire_425));
  TC_Or # (.UUID(64'd3711394974785431679 ^ UUID), .BIT_WIDTH(64'd8)) Or8_334 (.in0(wire_454), .in1(wire_193), .out(wire_226));
  TC_IndexerByte # (.UUID(64'd4264023620095411982 ^ UUID), .INDEX(64'd2)) IndexerByte_335 (.in(wire_130), .out(wire_454));
  TC_IndexerByte # (.UUID(64'd796235321624113339 ^ UUID), .INDEX(64'd3)) IndexerByte_336 (.in(wire_130), .out(wire_193));
  TC_Or # (.UUID(64'd327732458594941209 ^ UUID), .BIT_WIDTH(64'd8)) Or8_337 (.in0(wire_295), .in1(wire_384), .out(wire_342));
  TC_IndexerByte # (.UUID(64'd3956712446924886094 ^ UUID), .INDEX(64'd0)) IndexerByte_338 (.in(wire_130), .out(wire_295));
  TC_IndexerByte # (.UUID(64'd1400772416136704303 ^ UUID), .INDEX(64'd1)) IndexerByte_339 (.in(wire_130), .out(wire_384));
  TC_IndexerBit # (.UUID(64'd1173845344013116050 ^ UUID), .INDEX(64'd1)) IndexerBit_340 (.in({{56{1'b0}}, wire_196 }), .out(wire_408));
  TC_IndexerBit # (.UUID(64'd1993322735036255251 ^ UUID), .INDEX(64'd0)) IndexerBit_341 (.in({{56{1'b0}}, wire_196 }), .out(wire_400));
  TC_IndexerByte # (.UUID(64'd3961277922247604575 ^ UUID), .INDEX(64'd1)) IndexerByte_342 (.in({{48{1'b0}}, wire_161 }), .out(wire_196));
  TC_Equal # (.UUID(64'd2356628521336734568 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_343 (.in0(wire_256), .in1(wire_360), .out(wire_189));
  TC_Decoder3 # (.UUID(64'd1801936883088569704 ^ UUID)) Decoder3_344 (.dis(1'd0), .sel0(wire_401), .sel1(wire_375), .sel2(wire_115), .out0(), .out1(wire_4), .out2(wire_53), .out3(wire_223), .out4(wire_70), .out5(wire_101), .out6(wire_234), .out7(wire_411));
  TC_Constant # (.UUID(64'd1585905313389045148 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hC)) Constant8_345 (.out(wire_158));
  TC_Constant # (.UUID(64'd2027111329008812144 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hF)) Constant8_346 (.out(wire_473));
  TC_Switch # (.UUID(64'd510551550864988543 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_347 (.en(wire_223), .in(wire_473), .out(wire_168_2));
  TC_Switch # (.UUID(64'd4502977694884899110 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_348 (.en(wire_70), .in(wire_321), .out(wire_168_3));
  TC_Switch # (.UUID(64'd3444062419586535966 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_349 (.en(wire_101), .in(wire_388), .out(wire_168_4));
  TC_Switch # (.UUID(64'd3183065406337993090 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_350 (.en(wire_234), .in(wire_458), .out(wire_168_5));
  TC_Switch # (.UUID(64'd1881773228960447456 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_351 (.en(wire_411), .in(wire_210), .out(wire_168_6));
  TC_Constant # (.UUID(64'd287901269017399935 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h3)) Constant8_352 (.out(wire_465));
  TC_Not # (.UUID(64'd4058720228885546351 ^ UUID), .BIT_WIDTH(64'd1)) Not_353 (.in(wire_110), .out(wire_96));
  TC_Not # (.UUID(64'd781355532887995363 ^ UUID), .BIT_WIDTH(64'd1)) Not_354 (.in(wire_89), .out(wire_376));
  TC_Constant # (.UUID(64'd1765915980830865190 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h30)) Constant8_355 (.out(wire_321));
  TC_Switch # (.UUID(64'd4225563134404076393 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_356 (.en(wire_121), .in(wire_275), .out(wire_247));
  TC_IndexerBit # (.UUID(64'd1789832590864253294 ^ UUID), .INDEX(64'd7)) IndexerBit_357 (.in({{56{1'b0}}, wire_71 }), .out(wire_401));
  TC_IndexerBit # (.UUID(64'd423971802287147989 ^ UUID), .INDEX(64'd6)) IndexerBit_358 (.in({{56{1'b0}}, wire_71 }), .out(wire_375));
  TC_IndexerBit # (.UUID(64'd1849277145339495488 ^ UUID), .INDEX(64'd5)) IndexerBit_359 (.in({{56{1'b0}}, wire_71 }), .out(wire_115));
  TC_IndexerBit # (.UUID(64'd4348519509755259029 ^ UUID), .INDEX(64'd3)) IndexerBit_360 (.in({{56{1'b0}}, wire_71 }), .out(wire_59));
  TC_Switch # (.UUID(64'd139048722458446562 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_361 (.en(wire_53), .in(wire_158), .out(wire_168_1));
  TC_Switch # (.UUID(64'd1697328634740595572 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_362 (.en(wire_4), .in(wire_465), .out(wire_168_0));
  TC_Constant # (.UUID(64'd1476689218459702448 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h33)) Constant8_363 (.out(wire_388));
  TC_Constant # (.UUID(64'd3379970477126171844 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h3C)) Constant8_364 (.out(wire_458));
  TC_Constant # (.UUID(64'd304614014913386600 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h3F)) Constant8_365 (.out(wire_210));
  TC_Splitter16 # (.UUID(64'd3188721477555287760 ^ UUID)) Splitter16_366 (.in(wire_84[15:0]), .out0(), .out1(wire_256));
  TC_IndexerBit # (.UUID(64'd4049253696932042587 ^ UUID), .INDEX(64'd4)) IndexerBit_367 (.in({{56{1'b0}}, wire_71 }), .out(wire_54));
  TC_IndexerBit # (.UUID(64'd2814082116448811773 ^ UUID), .INDEX(64'd0)) IndexerBit_368 (.in({{48{1'b0}}, wire_161 }), .out(wire_10));
  TC_IndexerBit # (.UUID(64'd614485199549654646 ^ UUID), .INDEX(64'd1)) IndexerBit_369 (.in({{48{1'b0}}, wire_161 }), .out(wire_86));
  TC_IndexerBit # (.UUID(64'd3555852759017918092 ^ UUID), .INDEX(64'd2)) IndexerBit_370 (.in({{48{1'b0}}, wire_161 }), .out(wire_396));
  TC_IndexerBit # (.UUID(64'd1209262827994864386 ^ UUID), .INDEX(64'd3)) IndexerBit_371 (.in({{48{1'b0}}, wire_161 }), .out(wire_121));
  TC_Program # (.UUID(64'd3721980137216604240 ^ UUID), .WORD_WIDTH(64'd8), .DEFAULT_FILE_NAME("Program_33A7213703DAF850.w8.bin"), .ARG_SIG("Program_33A7213703DAF850=%s")) Program_372 (.clk(clk), .rst(rst), .address(wire_5), .out0(wire_156), .out1(), .out2(), .out3());
  TC_Splitter16 # (.UUID(64'd4461787469973933422 ^ UUID)) Splitter16_373 (.in(wire_84[15:0]), .out0(), .out1(wire_441));
  TC_Equal # (.UUID(64'd1988770091565985332 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_374 (.in0(wire_441), .in1(wire_102), .out(wire_385));
  TC_Constant # (.UUID(64'd2565543928344869306 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h5)) Constant8_375 (.out(wire_102));
  TC_Switch # (.UUID(64'd4105771623231641306 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_376 (.en(wire_385), .in(wire_156[15:0]), .out(wire_15_19[15:0]));
  TC_Equal # (.UUID(64'd551722571517782638 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_377 (.in0(16'd0), .in1(wire_6), .out(wire_106));
  TC_Or # (.UUID(64'd611236309732699826 ^ UUID), .BIT_WIDTH(64'd32)) Or32_378 (.in0({{31{1'b0}}, wire_328 }), .in1(wire_3), .out(wire_45));
  TC_DotMatrixDisplay # (.UUID(64'd1738323329834897739 ^ UUID)) DotMatrixDisplay_379 (.clk(clk), .rst(rst), .en_y(wire_45[0:0]), .en_x(wire_139[0:0]), .color_info(wire_45), .pixel_info(wire_139));
  TC_DotMatrixDisplay # (.UUID(64'd4354289896240283042 ^ UUID)) DotMatrixDisplay_380 (.clk(clk), .rst(rst), .en_y(wire_27[0:0]), .en_x(wire_139[0:0]), .color_info(wire_27), .pixel_info(wire_139));
  TC_Register # (.UUID(64'd4364107987795409853 ^ UUID), .BIT_WIDTH(64'd16)) Register16_381 (.clk(clk), .rst(rst), .load(wire_138), .save(wire_138), .in(wire_105), .out(wire_190));
  TC_Constant # (.UUID(64'd1415884859697557611 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_382 (.out(wire_37));
  TC_IndexerBit # (.UUID(64'd535377880148297947 ^ UUID), .INDEX(64'd3)) IndexerBit_383 (.in({{56{1'b0}}, wire_163 }), .out(wire_114));
  TC_Register # (.UUID(64'd2160598746671012754 ^ UUID), .BIT_WIDTH(64'd16)) Register16_384 (.clk(clk), .rst(rst), .load(wire_32), .save(wire_32), .in(wire_273), .out(wire_46));
  TC_Add # (.UUID(64'd1442806402229030427 ^ UUID), .BIT_WIDTH(64'd16)) Add16_385 (.in0(wire_132), .in1(wire_382), .ci(1'd0), .out(wire_73), .co());
  TC_Or # (.UUID(64'd2188959817660993009 ^ UUID), .BIT_WIDTH(64'd1)) Or_386 (.in0(wire_23), .in1(wire_66), .out(wire_32));
  TC_IndexerBit # (.UUID(64'd3588176080026118662 ^ UUID), .INDEX(64'd2)) IndexerBit_387 (.in({{56{1'b0}}, wire_163 }), .out(wire_289));
  TC_Mux # (.UUID(64'd4063471477342436371 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_388 (.sel(wire_66), .in0(wire_309), .in1(wire_46), .out(wire_132));
  TC_Mux # (.UUID(64'd527759690959107192 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_389 (.sel(wire_114), .in0(wire_165), .in1(wire_190), .out(wire_280));
  TC_Switch # (.UUID(64'd1362725833065582892 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_390 (.en(wire_289), .in(wire_105), .out(wire_165));
  TC_Switch # (.UUID(64'd1756831740426205013 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_391 (.en(wire_23), .in(wire_273), .out(wire_309));
  TC_Add # (.UUID(64'd2930665708224337659 ^ UUID), .BIT_WIDTH(64'd16)) Add16_392 (.in0(wire_190), .in1(wire_291), .ci(1'd0), .out(wire_105), .co());
  TC_Constant # (.UUID(64'd3137150186803814383 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hF0)) Constant8_393 (.out(wire_420));
  TC_Add # (.UUID(64'd432537638553101254 ^ UUID), .BIT_WIDTH(64'd16)) Add16_394 (.in0(wire_46), .in1(wire_413), .ci(1'd0), .out(wire_273), .co());
  TC_IndexerBit # (.UUID(64'd561707948535025464 ^ UUID), .INDEX(64'd4)) IndexerBit_395 (.in({{56{1'b0}}, wire_163 }), .out(wire_464));
  TC_Constant # (.UUID(64'd1695694096694981758 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_396 (.out(wire_173));
  TC_IndexerBit # (.UUID(64'd2331812482237933900 ^ UUID), .INDEX(64'd0)) IndexerBit_397 (.in({{56{1'b0}}, wire_149 }), .out(wire_359));
  TC_Neg # (.UUID(64'd1821476619534246961 ^ UUID), .BIT_WIDTH(64'd16)) Neg16_398 (.in({{8{1'b0}}, wire_173 }), .out(wire_63));
  TC_Mux # (.UUID(64'd1539425850473868597 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_399 (.sel(wire_464), .in0(wire_63), .in1({{8{1'b0}}, wire_173 }), .out(wire_413));
  TC_Mux # (.UUID(64'd3572805427243657698 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_400 (.sel(wire_289), .in0(wire_405), .in1({{8{1'b0}}, wire_37 }), .out(wire_291));
  TC_Neg # (.UUID(64'd2090057048615449572 ^ UUID), .BIT_WIDTH(64'd16)) Neg16_401 (.in({{8{1'b0}}, wire_37 }), .out(wire_405));
  TC_Constant # (.UUID(64'd245854699811937909 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h4)) Constant8_402 (.out(wire_360));
  TC_Splitter16 # (.UUID(64'd2039892175404791041 ^ UUID)) Splitter16_403 (.in(wire_255), .out0(wire_44), .out1(wire_230));
  TC_Constant # (.UUID(64'd886114160304713632 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hF8)) Constant8_404 (.out(wire_217));
  TC_And # (.UUID(64'd3416275225866990928 ^ UUID), .BIT_WIDTH(64'd8)) And8_405 (.in0(wire_217), .in1(wire_230), .out(wire_71));
  TC_Maker16 # (.UUID(64'd3199117322193596026 ^ UUID)) Maker16_406 (.in0(wire_209), .in1(wire_335), .out(wire_161));
  TC_Shr # (.UUID(64'd3593779976046315825 ^ UUID), .BIT_WIDTH(64'd8)) Shr8_407 (.in(wire_402), .shift(wire_208), .out(wire_335));
  TC_Switch # (.UUID(64'd4048603805359796154 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_408 (.en(wire_189), .in(wire_5), .out(wire_255));
  TC_Mul # (.UUID(64'd2182290031091560800 ^ UUID), .BIT_WIDTH(64'd8)) Mul8_409 (.in0(wire_251), .in1(wire_468), .out0(wire_55), .out1());
  TC_Constant # (.UUID(64'd3702906280545993063 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h8)) Constant8_410 (.out(wire_251));
  TC_Constant # (.UUID(64'd182979028355080598 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6)) Constant8_411 (.out(wire_235));
  TC_Mul # (.UUID(64'd65965927015369652 ^ UUID), .BIT_WIDTH(64'd8)) DivMod8_412 (.in0(wire_203[7:0]), .in1(wire_235), .out0(wire_209), .out1(wire_468));
  TC_Constant # (.UUID(64'd1209373824649557251 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h5)) Constant8_413 (.out(wire_423));
  TC_And # (.UUID(64'd3192677659232933832 ^ UUID), .BIT_WIDTH(64'd8)) And8_414 (.in0(wire_230), .in1(wire_358), .out(wire_447));
  TC_Constant # (.UUID(64'd3278513372338526303 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7)) Constant8_415 (.out(wire_326));
  TC_And # (.UUID(64'd333727324415720762 ^ UUID), .BIT_WIDTH(64'd8)) And8_416 (.in0(wire_402), .in1(wire_326), .out(wire_288));
  TC_Add # (.UUID(64'd3323828643250169126 ^ UUID), .BIT_WIDTH(64'd8)) Add8_417 (.in0(wire_55), .in1(wire_288), .ci(1'd0), .out(wire_249), .co());
  TC_Maker16 # (.UUID(64'd4018174165342853046 ^ UUID)) Maker16_418 (.in0(wire_44), .in1(wire_447), .out(wire_348));
  TC_And # (.UUID(64'd3586445645766121843 ^ UUID), .BIT_WIDTH(64'd8)) And8_419 (.in0(wire_44), .in1(wire_337), .out(wire_402));
  TC_Shr # (.UUID(64'd700522554472714991 ^ UUID), .BIT_WIDTH(64'd16)) Shr16_420 (.in(wire_348), .shift(wire_423), .out(wire_203));
  TC_Constant # (.UUID(64'd826175156228145649 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1F)) Constant8_421 (.out(wire_337));
  TC_Constant # (.UUID(64'd1842362314523162062 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7)) Constant8_422 (.out(wire_358));
  TC_Constant # (.UUID(64'd811789851201528647 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h3)) Constant8_423 (.out(wire_208));
  TC_IOSwitch # (.UUID(64'd2846053541171193881 ^ UUID), .BIT_WIDTH(64'd8)) LevelOutputArch_424 (.in(wire_5[7:0]), .en(wire_319), .out(arch_output_value));
  TC_Switch # (.UUID(64'd210661621448949326 ^ UUID), .BIT_WIDTH(64'd8)) LevelInputArch_425 (.en(wire_151), .in(arch_input_value), .out(wire_15_20[7:0]));
  TC_Splitter16 # (.UUID(64'd2775342692045340835 ^ UUID)) Splitter16_426 (.in(wire_84[15:0]), .out0(), .out1(wire_306));
  TC_Equal # (.UUID(64'd4532639728004948159 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_427 (.in0(wire_306), .in1(wire_199), .out(wire_264));
  TC_Equal # (.UUID(64'd3745587913460272427 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_428 (.in0(wire_322), .in1(wire_306), .out(wire_415));
  TC_Constant # (.UUID(64'd951998662890801082 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6)) Constant8_429 (.out(wire_322));
  TC_Constant # (.UUID(64'd2262634952183580731 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7)) Constant8_430 (.out(wire_199));
  TC_Switch # (.UUID(64'd1419008802292368204 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_431 (.en(wire_25), .in(wire_415), .out(wire_151));
  TC_Clock # (.UUID(64'd150335021447124340 ^ UUID)) Clock_432 (.clk(clk), .rst(rst), .out(wire_25));
  TC_Switch # (.UUID(64'd3781955660154943019 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_433 (.en(wire_277), .in(wire_264), .out(wire_319));
  TC_Not # (.UUID(64'd248590985388437467 ^ UUID), .BIT_WIDTH(64'd1)) Not_434 (.in(wire_25), .out(wire_277));
  TC_RamDualLoad # (.UUID(64'd1162091816344660036 ^ UUID), .WORD_WIDTH(64'd16), .WORD_COUNT(64'd65536)) RamDualLoad_435 (.clk(clk), .rst(rst), .load0(wire_74), .save(wire_451), .address0({{16{1'b0}}, wire_143 }), .in({{48{1'b0}}, wire_177 }), .load1(wire_28), .address1({{16{1'b0}}, wire_227 }), .out0(wire_38), .out1(wire_315));
  TC_Ram # (.UUID(64'd2071862132571227302 ^ UUID), .WORD_WIDTH(64'd16), .WORD_COUNT(64'd65536)) Ram_436 (.clk(clk), .rst(rst), .load(wire_106), .save(wire_131), .address({{16{1'b0}}, wire_13 }), .in0({{48{1'b0}}, wire_6 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_343), .out1(), .out2(), .out3());
  TC_FileLoader # (.UUID(64'd1149854990232492044 ^ UUID), .DEFAULT_FILE_NAME("test.dat")) FileLoader_437 (.clk(clk), .rst(rst), .en(wire_48), .address({{48{1'b0}}, wire_5 }), .out(wire_15_13));
  TC_Splitter16 # (.UUID(64'd2684349980131024015 ^ UUID)) Splitter16_438 (.in(wire_84[15:0]), .out0(), .out1(wire_353));
  TC_Equal # (.UUID(64'd4369488988257915881 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_439 (.in0(wire_353), .in1(wire_344), .out(wire_48));
  TC_Constant # (.UUID(64'd3823619217162964047 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7)) Constant8_440 (.out(wire_344));
  TC_Ror # (.UUID(64'd445352019034615982 ^ UUID), .BIT_WIDTH(64'd16)) Ror16_441 (.in(wire_5), .shift(wire_24[7:0]), .out(wire_455));
  TC_IndexerBit # (.UUID(64'd815489067524461103 ^ UUID), .INDEX(64'd6)) IndexerBit_442 (.in({{56{1'b0}}, wire_249 }), .out(wire_91));

  wire [0:0] wire_0;
  wire [0:0] wire_1;
  wire [0:0] wire_2;
  wire [0:0] wire_2_0;
  wire [0:0] wire_2_1;
  wire [0:0] wire_2_2;
  wire [0:0] wire_2_3;
  wire [0:0] wire_2_4;
  wire [0:0] wire_2_5;
  wire [0:0] wire_2_6;
  wire [0:0] wire_2_7;
  wire [0:0] wire_2_8;
  wire [0:0] wire_2_9;
  assign wire_2 = wire_2_0|wire_2_1|wire_2_2|wire_2_3|wire_2_4|wire_2_5|wire_2_6|wire_2_7|wire_2_8|wire_2_9;
  wire [31:0] wire_3;
  wire [0:0] wire_4;
  wire [15:0] wire_5;
  wire [15:0] wire_5_0;
  wire [15:0] wire_5_1;
  assign wire_5 = wire_5_0|wire_5_1;
  wire [15:0] wire_6;
  wire [0:0] wire_7;
  wire [7:0] wire_8;
  wire [31:0] wire_9;
  wire [0:0] wire_10;
  wire [63:0] wire_11;
  wire [0:0] wire_12;
  wire [15:0] wire_13;
  wire [0:0] wire_14;
  wire [63:0] wire_15;
  wire [63:0] wire_15_0;
  wire [63:0] wire_15_1;
  wire [63:0] wire_15_2;
  wire [63:0] wire_15_3;
  wire [63:0] wire_15_4;
  wire [63:0] wire_15_5;
  wire [63:0] wire_15_6;
  wire [63:0] wire_15_7;
  wire [63:0] wire_15_8;
  wire [63:0] wire_15_9;
  wire [63:0] wire_15_10;
  wire [63:0] wire_15_11;
  wire [63:0] wire_15_12;
  wire [63:0] wire_15_13;
  wire [63:0] wire_15_14;
  wire [63:0] wire_15_15;
  wire [63:0] wire_15_16;
  wire [63:0] wire_15_17;
  wire [63:0] wire_15_18;
  wire [63:0] wire_15_19;
  wire [63:0] wire_15_20;
  assign wire_15 = wire_15_0|wire_15_1|wire_15_2|wire_15_3|wire_15_4|wire_15_5|wire_15_6|wire_15_7|wire_15_8|wire_15_9|wire_15_10|wire_15_11|wire_15_12|wire_15_13|wire_15_14|wire_15_15|wire_15_16|wire_15_17|wire_15_18|wire_15_19|wire_15_20;
  wire [0:0] wire_16;
  wire [15:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [15:0] wire_21;
  wire [15:0] wire_21_0;
  wire [15:0] wire_21_1;
  wire [15:0] wire_21_2;
  assign wire_21 = wire_21_0|wire_21_1|wire_21_2;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [15:0] wire_24;
  wire [15:0] wire_24_0;
  wire [15:0] wire_24_1;
  assign wire_24 = wire_24_0|wire_24_1;
  wire [0:0] wire_25;
  wire [63:0] wire_26;
  wire [31:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  assign wire_34 = 0;
  wire [0:0] wire_35;
  wire [15:0] wire_36;
  wire [7:0] wire_37;
  wire [63:0] wire_38;
  wire [0:0] wire_39;
  wire [0:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [7:0] wire_44;
  wire [31:0] wire_45;
  wire [15:0] wire_46;
  wire [15:0] wire_47;
  wire [0:0] wire_48;
  wire [0:0] wire_49;
  wire [31:0] wire_50;
  wire [0:0] wire_51;
  wire [15:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  wire [7:0] wire_55;
  wire [0:0] wire_56;
  wire [15:0] wire_57;
  wire [15:0] wire_58;
  wire [0:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [31:0] wire_62;
  wire [15:0] wire_63;
  wire [0:0] wire_64;
  wire [7:0] wire_65;
  wire [0:0] wire_66;
  wire [0:0] wire_67;
  wire [31:0] wire_68;
  wire [0:0] wire_69;
  wire [0:0] wire_70;
  wire [7:0] wire_71;
  wire [0:0] wire_72;
  wire [15:0] wire_73;
  wire [0:0] wire_74;
  wire [0:0] wire_75;
  wire [0:0] wire_76;
  wire [0:0] wire_77;
  wire [0:0] wire_78;
  wire [0:0] wire_79;
  wire [0:0] wire_80;
  wire [0:0] wire_81;
  wire [63:0] wire_82;
  wire [0:0] wire_83;
  wire [63:0] wire_84;
  wire [0:0] wire_85;
  wire [0:0] wire_86;
  wire [0:0] wire_87;
  wire [15:0] wire_88;
  wire [0:0] wire_89;
  wire [0:0] wire_90;
  wire [0:0] wire_91;
  wire [15:0] wire_92;
  wire [0:0] wire_93;
  wire [0:0] wire_94;
  wire [0:0] wire_95;
  wire [0:0] wire_96;
  wire [15:0] wire_97;
  wire [15:0] wire_97_0;
  wire [15:0] wire_97_1;
  assign wire_97 = wire_97_0|wire_97_1;
  wire [31:0] wire_98;
  wire [7:0] wire_99;
  wire [0:0] wire_100;
  wire [0:0] wire_101;
  wire [7:0] wire_102;
  wire [0:0] wire_103;
  wire [15:0] wire_104;
  wire [15:0] wire_105;
  wire [0:0] wire_106;
  wire [0:0] wire_107;
  wire [0:0] wire_108;
  wire [0:0] wire_109;
  wire [0:0] wire_110;
  wire [63:0] wire_111;
  wire [15:0] wire_112;
  wire [63:0] wire_113;
  wire [0:0] wire_114;
  wire [0:0] wire_115;
  wire [0:0] wire_116;
  wire [31:0] wire_117;
  wire [15:0] wire_118;
  wire [0:0] wire_119;
  wire [0:0] wire_120;
  wire [0:0] wire_121;
  wire [0:0] wire_122;
  wire [0:0] wire_123;
  wire [15:0] wire_124;
  wire [15:0] wire_125;
  wire [0:0] wire_126;
  wire [0:0] wire_127;
  wire [15:0] wire_128;
  wire [31:0] wire_129;
  wire [63:0] wire_130;
  wire [0:0] wire_131;
  wire [15:0] wire_132;
  wire [31:0] wire_133;
  wire [0:0] wire_134;
  wire [31:0] wire_135;
  wire [0:0] wire_136;
  wire [15:0] wire_137;
  wire [0:0] wire_138;
  wire [63:0] wire_139;
  wire [63:0] wire_140;
  wire [0:0] wire_141;
  wire [63:0] wire_142;
  wire [15:0] wire_143;
  wire [15:0] wire_143_0;
  wire [15:0] wire_143_1;
  assign wire_143 = wire_143_0|wire_143_1;
  wire [0:0] wire_144;
  wire [0:0] wire_145;
  wire [0:0] wire_146;
  wire [15:0] wire_147;
  wire [0:0] wire_148;
  wire [7:0] wire_149;
  wire [0:0] wire_150;
  wire [0:0] wire_151;
  assign arch_input_enable = wire_151;
  wire [15:0] wire_152;
  wire [7:0] wire_153;
  wire [0:0] wire_154;
  wire [7:0] wire_155;
  wire [63:0] wire_156;
  wire [7:0] wire_157;
  wire [7:0] wire_158;
  wire [0:0] wire_159;
  wire [7:0] wire_160;
  wire [15:0] wire_161;
  wire [0:0] wire_162;
  wire [7:0] wire_163;
  wire [0:0] wire_164;
  wire [15:0] wire_165;
  wire [0:0] wire_166;
  wire [0:0] wire_167;
  wire [7:0] wire_168;
  wire [7:0] wire_168_0;
  wire [7:0] wire_168_1;
  wire [7:0] wire_168_2;
  wire [7:0] wire_168_3;
  wire [7:0] wire_168_4;
  wire [7:0] wire_168_5;
  wire [7:0] wire_168_6;
  assign wire_168 = wire_168_0|wire_168_1|wire_168_2|wire_168_3|wire_168_4|wire_168_5|wire_168_6;
  wire [0:0] wire_169;
  wire [0:0] wire_170;
  wire [0:0] wire_171;
  wire [0:0] wire_172;
  wire [7:0] wire_173;
  wire [15:0] wire_174;
  wire [0:0] wire_175;
  wire [0:0] wire_176;
  wire [15:0] wire_177;
  wire [0:0] wire_178;
  wire [0:0] wire_178_0;
  wire [0:0] wire_178_1;
  wire [0:0] wire_178_2;
  assign wire_178 = wire_178_0|wire_178_1|wire_178_2;
  wire [0:0] wire_179;
  wire [0:0] wire_180;
  wire [0:0] wire_181;
  wire [0:0] wire_182;
  wire [0:0] wire_183;
  wire [0:0] wire_184;
  wire [0:0] wire_185;
  wire [15:0] wire_186;
  wire [63:0] wire_187;
  wire [0:0] wire_188;
  wire [0:0] wire_189;
  wire [15:0] wire_190;
  wire [0:0] wire_191;
  wire [7:0] wire_192;
  wire [7:0] wire_193;
  wire [0:0] wire_194;
  wire [7:0] wire_195;
  wire [7:0] wire_196;
  wire [7:0] wire_197;
  wire [0:0] wire_198;
  wire [7:0] wire_199;
  wire [0:0] wire_200;
  wire [0:0] wire_201;
  wire [0:0] wire_202;
  wire [15:0] wire_203;
  wire [0:0] wire_204;
  wire [7:0] wire_205;
  wire [0:0] wire_206;
  wire [0:0] wire_207;
  wire [7:0] wire_208;
  wire [7:0] wire_209;
  wire [7:0] wire_210;
  wire [0:0] wire_211;
  wire [0:0] wire_212;
  wire [0:0] wire_213;
  wire [7:0] wire_214;
  wire [0:0] wire_215;
  wire [0:0] wire_216;
  wire [7:0] wire_217;
  wire [0:0] wire_218;
  wire [15:0] wire_219;
  wire [0:0] wire_220;
  wire [0:0] wire_221;
  wire [0:0] wire_222;
  wire [0:0] wire_223;
  wire [7:0] wire_224;
  wire [63:0] wire_225;
  wire [7:0] wire_226;
  wire [15:0] wire_227;
  wire [0:0] wire_228;
  wire [15:0] wire_229;
  wire [7:0] wire_230;
  wire [31:0] wire_231;
  wire [0:0] wire_232;
  wire [0:0] wire_233;
  wire [0:0] wire_234;
  wire [7:0] wire_235;
  wire [0:0] wire_236;
  wire [15:0] wire_237;
  wire [0:0] wire_238;
  wire [0:0] wire_239;
  wire [0:0] wire_240;
  wire [0:0] wire_241;
  wire [0:0] wire_242;
  wire [15:0] wire_243;
  wire [0:0] wire_244;
  wire [0:0] wire_245;
  wire [0:0] wire_246;
  wire [0:0] wire_247;
  wire [31:0] wire_248;
  wire [7:0] wire_249;
  wire [0:0] wire_250;
  wire [7:0] wire_251;
  wire [7:0] wire_252;
  wire [0:0] wire_253;
  wire [7:0] wire_254;
  wire [15:0] wire_255;
  wire [7:0] wire_256;
  wire [15:0] wire_257;
  wire [0:0] wire_258;
  wire [7:0] wire_259;
  wire [0:0] wire_260;
  wire [7:0] wire_261;
  wire [7:0] wire_262;
  wire [0:0] wire_263;
  wire [0:0] wire_264;
  wire [0:0] wire_265;
  wire [0:0] wire_266;
  wire [0:0] wire_267;
  wire [0:0] wire_268;
  wire [0:0] wire_269;
  wire [0:0] wire_270;
  wire [0:0] wire_271;
  wire [0:0] wire_272;
  wire [15:0] wire_273;
  wire [0:0] wire_274;
  wire [0:0] wire_275;
  wire [0:0] wire_276;
  wire [0:0] wire_277;
  wire [0:0] wire_278;
  wire [0:0] wire_279;
  wire [15:0] wire_280;
  wire [0:0] wire_281;
  wire [15:0] wire_282;
  wire [0:0] wire_283;
  wire [0:0] wire_284;
  wire [0:0] wire_285;
  wire [0:0] wire_286;
  wire [0:0] wire_287;
  wire [7:0] wire_288;
  wire [0:0] wire_289;
  wire [15:0] wire_290;
  wire [15:0] wire_291;
  wire [0:0] wire_292;
  wire [63:0] wire_293;
  wire [0:0] wire_294;
  wire [7:0] wire_295;
  wire [0:0] wire_296;
  wire [0:0] wire_297;
  wire [0:0] wire_298;
  wire [7:0] wire_299;
  wire [0:0] wire_300;
  wire [0:0] wire_301;
  wire [0:0] wire_302;
  wire [0:0] wire_303;
  wire [7:0] wire_304;
  wire [0:0] wire_305;
  wire [7:0] wire_306;
  wire [0:0] wire_307;
  wire [0:0] wire_308;
  wire [15:0] wire_309;
  wire [0:0] wire_310;
  wire [0:0] wire_311;
  wire [0:0] wire_312;
  wire [0:0] wire_313;
  wire [0:0] wire_314;
  wire [63:0] wire_315;
  wire [0:0] wire_316;
  wire [0:0] wire_317;
  wire [63:0] wire_318;
  wire [0:0] wire_319;
  assign arch_output_enable = wire_319;
  wire [0:0] wire_320;
  wire [7:0] wire_321;
  wire [7:0] wire_322;
  wire [7:0] wire_323;
  wire [0:0] wire_324;
  wire [0:0] wire_325;
  wire [7:0] wire_326;
  wire [63:0] wire_327;
  wire [0:0] wire_328;
  wire [0:0] wire_329;
  wire [0:0] wire_330;
  wire [0:0] wire_331;
  wire [7:0] wire_332;
  wire [63:0] wire_333;
  wire [0:0] wire_334;
  wire [7:0] wire_335;
  wire [15:0] wire_336;
  wire [7:0] wire_337;
  wire [0:0] wire_338;
  wire [0:0] wire_339;
  wire [7:0] wire_340;
  wire [0:0] wire_341;
  wire [7:0] wire_342;
  wire [63:0] wire_343;
  wire [7:0] wire_344;
  wire [7:0] wire_345;
  wire [0:0] wire_346;
  wire [0:0] wire_347;
  wire [15:0] wire_348;
  wire [0:0] wire_349;
  wire [7:0] wire_350;
  wire [0:0] wire_351;
  wire [7:0] wire_352;
  wire [7:0] wire_353;
  wire [0:0] wire_354;
  wire [0:0] wire_355;
  wire [7:0] wire_356;
  wire [15:0] wire_357;
  wire [7:0] wire_358;
  wire [0:0] wire_359;
  wire [7:0] wire_360;
  wire [0:0] wire_361;
  wire [0:0] wire_362;
  wire [0:0] wire_363;
  wire [0:0] wire_364;
  wire [0:0] wire_365;
  wire [0:0] wire_366;
  wire [7:0] wire_367;
  wire [0:0] wire_368;
  wire [7:0] wire_369;
  wire [0:0] wire_370;
  wire [7:0] wire_371;
  wire [0:0] wire_372;
  wire [15:0] wire_373;
  wire [7:0] wire_374;
  wire [0:0] wire_375;
  wire [0:0] wire_376;
  wire [0:0] wire_377;
  wire [0:0] wire_378;
  wire [0:0] wire_379;
  wire [0:0] wire_380;
  wire [7:0] wire_381;
  wire [15:0] wire_382;
  wire [0:0] wire_383;
  wire [7:0] wire_384;
  wire [0:0] wire_385;
  wire [15:0] wire_386;
  wire [15:0] wire_387;
  wire [7:0] wire_388;
  wire [0:0] wire_389;
  wire [15:0] wire_390;
  wire [0:0] wire_391;
  wire [15:0] wire_392;
  wire [0:0] wire_393;
  wire [0:0] wire_394;
  wire [0:0] wire_395;
  wire [0:0] wire_396;
  wire [0:0] wire_397;
  wire [0:0] wire_398;
  wire [0:0] wire_399;
  wire [0:0] wire_400;
  wire [0:0] wire_401;
  wire [7:0] wire_402;
  wire [7:0] wire_403;
  wire [7:0] wire_404;
  wire [15:0] wire_405;
  wire [0:0] wire_406;
  wire [15:0] wire_407;
  wire [0:0] wire_408;
  wire [0:0] wire_409;
  wire [0:0] wire_410;
  wire [0:0] wire_411;
  wire [7:0] wire_412;
  wire [15:0] wire_413;
  wire [63:0] wire_414;
  wire [0:0] wire_415;
  wire [0:0] wire_416;
  wire [0:0] wire_417;
  wire [0:0] wire_418;
  wire [0:0] wire_419;
  wire [7:0] wire_420;
  wire [7:0] wire_421;
  wire [0:0] wire_422;
  wire [7:0] wire_423;
  wire [7:0] wire_424;
  wire [7:0] wire_425;
  wire [0:0] wire_426;
  wire [0:0] wire_427;
  wire [7:0] wire_428;
  wire [0:0] wire_429;
  wire [0:0] wire_430;
  wire [0:0] wire_431;
  wire [0:0] wire_432;
  wire [15:0] wire_433;
  wire [0:0] wire_434;
  wire [0:0] wire_435;
  wire [7:0] wire_436;
  wire [0:0] wire_437;
  wire [0:0] wire_438;
  wire [0:0] wire_439;
  wire [0:0] wire_440;
  wire [7:0] wire_441;
  wire [0:0] wire_442;
  wire [0:0] wire_443;
  wire [0:0] wire_444;
  wire [0:0] wire_445;
  wire [7:0] wire_446;
  wire [7:0] wire_447;
  wire [0:0] wire_448;
  wire [0:0] wire_449;
  wire [0:0] wire_450;
  wire [0:0] wire_451;
  wire [0:0] wire_452;
  wire [0:0] wire_453;
  wire [7:0] wire_454;
  wire [15:0] wire_455;
  wire [0:0] wire_456;
  wire [0:0] wire_457;
  wire [7:0] wire_458;
  wire [0:0] wire_459;
  wire [7:0] wire_460;
  wire [0:0] wire_461;
  wire [0:0] wire_462;
  wire [0:0] wire_463;
  wire [0:0] wire_464;
  wire [7:0] wire_465;
  wire [0:0] wire_466;
  wire [0:0] wire_467;
  wire [7:0] wire_468;
  wire [0:0] wire_469;
  wire [0:0] wire_470;
  wire [7:0] wire_471;
  wire [0:0] wire_472;
  wire [7:0] wire_473;
  wire [0:0] wire_474;
  wire [0:0] wire_475;
  wire [0:0] wire_476;

endmodule
