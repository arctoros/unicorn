module Unicornz_128x128 (clk, rst, arch_output_enable, arch_output_value, arch_input_enable, arch_input_value);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  output  wire [0:0] arch_output_enable;
  output  wire [7:0] arch_output_value;
  output  wire [0:0] arch_input_enable;
  input  wire [7:0] arch_input_value;

  TC_Program # (.UUID(64'd2054094413772625173 ^ UUID), .WORD_WIDTH(64'd16), .DEFAULT_FILE_NAME("Program_1C819BFC7C081515.w16.bin"), .ARG_SIG("Program_1C819BFC7C081515=%s")) Program_0 (.clk(clk), .rst(rst), .address(wire_55), .out0(wire_21), .out1(wire_104), .out2(wire_327), .out3(wire_424));
  TC_Decoder3 # (.UUID(64'd2564548179517358600 ^ UUID)) Decoder3_1 (.dis(wire_146), .sel0(wire_99), .sel1(wire_96), .sel2(wire_115), .out0(wire_473), .out1(wire_196), .out2(wire_492), .out3(wire_333), .out4(wire_252), .out5(wire_465), .out6(wire_418), .out7(wire_463));
  TC_Decoder3 # (.UUID(64'd3856915764158948127 ^ UUID)) Decoder3_2 (.dis(wire_226), .sel0(wire_99), .sel1(wire_96), .sel2(wire_115), .out0(wire_254), .out1(wire_456), .out2(wire_339), .out3(wire_495), .out4(wire_407), .out5(wire_156), .out6(wire_383), .out7(wire_453));
  TC_Decoder3 # (.UUID(64'd469263968959042607 ^ UUID)) Decoder3_3 (.dis(wire_396), .sel0(wire_99), .sel1(wire_96), .sel2(wire_115), .out0(wire_464), .out1(wire_378), .out2(wire_451), .out3(wire_408), .out4(wire_440), .out5(wire_432), .out6(wire_347), .out7(wire_356));
  TC_Decoder3 # (.UUID(64'd2355515313084503399 ^ UUID)) Decoder3_4 (.dis(wire_127), .sel0(wire_99), .sel1(wire_96), .sel2(wire_115), .out0(wire_372), .out1(wire_370), .out2(wire_455), .out3(wire_219), .out4(wire_260), .out5(wire_297), .out6(wire_350), .out7(wire_420));
  TC_Maker8 # (.UUID(64'd3412742270897961611 ^ UUID)) Maker8_5 (.in0(wire_473), .in1(wire_196), .in2(wire_492), .in3(wire_333), .in4(wire_252), .in5(wire_465), .in6(wire_418), .in7(wire_463), .out(wire_269));
  TC_Maker8 # (.UUID(64'd2545466735680713447 ^ UUID)) Maker8_6 (.in0(wire_254), .in1(wire_456), .in2(wire_339), .in3(wire_495), .in4(wire_407), .in5(wire_156), .in6(wire_383), .in7(wire_453), .out(wire_364));
  TC_Maker8 # (.UUID(64'd2498328128700172685 ^ UUID)) Maker8_7 (.in0(wire_464), .in1(wire_378), .in2(wire_451), .in3(wire_408), .in4(wire_440), .in5(wire_432), .in6(wire_347), .in7(wire_356), .out(wire_483));
  TC_Maker8 # (.UUID(64'd3307623088924666213 ^ UUID)) Maker8_8 (.in0(wire_372), .in1(wire_370), .in2(wire_455), .in3(wire_219), .in4(wire_260), .in5(wire_297), .in6(wire_350), .in7(wire_420), .out(wire_27));
  TC_Maker32 # (.UUID(64'd3223173008764962790 ^ UUID)) Maker32_9 (.in0(wire_27), .in1(wire_483), .in2(wire_364), .in3(wire_269), .out(wire_48));
  TC_Switch # (.UUID(64'd1126631217811470669 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_10 (.en(wire_295), .in(wire_50), .out(wire_155));
  TC_Switch # (.UUID(64'd383016835864160285 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_11 (.en(wire_307), .in(wire_187), .out(wire_12_0));
  TC_Switch # (.UUID(64'd3140243124393805415 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_12 (.en(wire_417), .in(wire_25), .out(wire_101));
  TC_Switch # (.UUID(64'd1581886471977480656 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_13 (.en(wire_373), .in(wire_25), .out(wire_51_1));
  TC_Switch # (.UUID(64'd2241249704231886051 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_14 (.en(wire_240), .in(wire_327[15:0]), .out(wire_187));
  TC_Switch # (.UUID(64'd4100643114395522594 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_15 (.en(wire_267), .in(wire_104[15:0]), .out(wire_50_2));
  TC_Switch # (.UUID(64'd8725165111331077 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_16 (.en(wire_34), .in(wire_327[15:0]), .out(wire_50_1));
  TC_Switch # (.UUID(64'd3499335185666676498 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_17 (.en(wire_240), .in(wire_424[15:0]), .out(wire_50_0));
  TC_And3 # (.UUID(64'd2537048141319315915 ^ UUID), .BIT_WIDTH(64'd1)) And3_18 (.in0(wire_5), .in1(wire_296), .in2(wire_191), .out(wire_75));
  TC_Program # (.UUID(64'd388994960009383908 ^ UUID), .WORD_WIDTH(64'd32), .DEFAULT_FILE_NAME("Program_565FCDAEAC6CFE4.w32.bin"), .ARG_SIG("Program_565FCDAEAC6CFE4=%s")) Program_19 (.clk(clk), .rst(rst), .address({{8{1'b0}}, wire_235 }), .out0(wire_36), .out1(), .out2(), .out3());
  TC_Not # (.UUID(64'd2992010998666944854 ^ UUID), .BIT_WIDTH(64'd1)) Not_20 (.in(wire_220), .out(wire_423));
  TC_Switch # (.UUID(64'd92717477479612822 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_21 (.en(wire_142), .in(wire_326), .out(wire_151));
  TC_Counter # (.UUID(64'd388538542796967315 ^ UUID), .BIT_WIDTH(64'd16), .count(16'd1)) Counter16_22 (.clk(clk), .rst(rst), .save(wire_220), .in(wire_177), .out(wire_290));
  TC_Counter # (.UUID(64'd3159443906265585347 ^ UUID), .BIT_WIDTH(64'd16), .count(16'd1)) Counter16_23 (.clk(clk), .rst(rst), .save(wire_435), .in(wire_177), .out(wire_10));
  TC_DelayLine # (.UUID(64'd1367561201104940128 ^ UUID), .BIT_WIDTH(64'd16)) DelayLine16_24 (.clk(clk), .rst(rst), .in(wire_83[15:0]), .out(wire_326));
  TC_Switch # (.UUID(64'd4093327232412684622 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_25 (.en(wire_220), .in(wire_10), .out(wire_79_1));
  TC_Switch # (.UUID(64'd3521663283135285715 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_26 (.en(wire_423), .in(wire_290), .out(wire_79_0));
  TC_Mux # (.UUID(64'd3040671060942591441 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_27 (.sel(wire_142), .in0(wire_79), .in1(wire_151), .out(wire_55));
  TC_DelayLine # (.UUID(64'd1970975974056862148 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_28 (.clk(clk), .rst(rst), .in(wire_90), .out(wire_142));
  TC_DelayLine # (.UUID(64'd4083747472069111906 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_29 (.clk(clk), .rst(rst), .in(wire_220), .out(wire_435));
  TC_Not # (.UUID(64'd2703499132143664233 ^ UUID), .BIT_WIDTH(64'd1)) Not_30 (.in(wire_435), .out(wire_220));
  TC_Not # (.UUID(64'd668729040907233308 ^ UUID), .BIT_WIDTH(64'd1)) Not_31 (.in(wire_115), .out(wire_159));
  TC_Not # (.UUID(64'd1492999759409908823 ^ UUID), .BIT_WIDTH(64'd1)) Not_32 (.in(wire_99), .out(wire_249));
  TC_And3 # (.UUID(64'd3485287916682882951 ^ UUID), .BIT_WIDTH(64'd1)) And3_33 (.in0(wire_159), .in1(wire_96), .in2(wire_249), .out(wire_191));
  TC_Switch # (.UUID(64'd1180978168546894742 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_34 (.en(wire_75), .in(wire_75), .out(wire_100_1));
  TC_Switch # (.UUID(64'd3723419762929890741 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_35 (.en(wire_34), .in(wire_34), .out(wire_100_0));
  TC_Switch # (.UUID(64'd2050768528734077835 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_36 (.en(wire_240), .in(wire_240), .out(wire_100_2));
  TC_Switch # (.UUID(64'd3057161046631511266 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_37 (.en(wire_255), .in(wire_255), .out(wire_34));
  TC_Decoder2 # (.UUID(64'd3508168605160458460 ^ UUID)) Decoder2_38 (.sel0(wire_131), .sel1(wire_93), .out0(), .out1(), .out2(wire_195), .out3(wire_255));
  TC_Not # (.UUID(64'd1768466669334456870 ^ UUID), .BIT_WIDTH(64'd1)) Not_39 (.in(wire_75), .out(wire_203));
  TC_Not # (.UUID(64'd3282289532960715218 ^ UUID), .BIT_WIDTH(64'd1)) Not_40 (.in(wire_18), .out(wire_226));
  TC_Not # (.UUID(64'd1327891776776277559 ^ UUID), .BIT_WIDTH(64'd1)) Not_41 (.in(wire_86), .out(wire_396));
  TC_Not # (.UUID(64'd1982359815710823425 ^ UUID), .BIT_WIDTH(64'd1)) Not_42 (.in(wire_60), .out(wire_127));
  TC_Decoder2 # (.UUID(64'd2605064451303635720 ^ UUID)) Decoder2_43 (.sel0(wire_296), .sel1(wire_5), .out0(wire_60), .out1(wire_86), .out2(wire_18), .out3(wire_481));
  TC_Add # (.UUID(64'd3313543325696297390 ^ UUID), .BIT_WIDTH(64'd16)) Add16_44 (.in0(wire_55), .in1(wire_36[15:0]), .ci(1'd0), .out(wire_177), .co());
  TC_IndexerBit # (.UUID(64'd2196806765189308211 ^ UUID), .INDEX(64'd1)) IndexerBit_45 (.in(wire_36), .out(wire_93));
  TC_IndexerBit # (.UUID(64'd737839460036088508 ^ UUID), .INDEX(64'd0)) IndexerBit_46 (.in(wire_36), .out(wire_131));
  TC_IndexerBit # (.UUID(64'd2903462054980356400 ^ UUID), .INDEX(64'd2)) IndexerBit_47 (.in(wire_36), .out(wire_240));
  TC_Splitter8 # (.UUID(64'd3910511016620535394 ^ UUID)) Splitter8_48 (.in(wire_450), .out0(wire_342), .out1(wire_132), .out2(wire_63), .out3(wire_161), .out4(wire_124), .out5(wire_305), .out6(wire_110), .out7(wire_218));
  TC_IndexerByte # (.UUID(64'd2436263972142084427 ^ UUID), .INDEX(64'd1)) IndexerByte_49 (.in({{32{1'b0}}, wire_48 }), .out(wire_450));
  TC_Switch # (.UUID(64'd607808644696146469 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_50 (.en(wire_342), .in(wire_390), .out(wire_83_10[15:0]));
  TC_Switch # (.UUID(64'd2632353714035774615 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_51 (.en(wire_132), .in(wire_288), .out(wire_83_12[15:0]));
  TC_Switch # (.UUID(64'd2222450423847071001 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_52 (.en(wire_63), .in(wire_106), .out(wire_83_14[15:0]));
  TC_Switch # (.UUID(64'd3314256307520299439 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_53 (.en(wire_161), .in(wire_353), .out(wire_83_16[15:0]));
  TC_Switch # (.UUID(64'd2595134878720988598 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_54 (.en(wire_124), .in(wire_76), .out(wire_83_17[15:0]));
  TC_Switch # (.UUID(64'd1299382207876995858 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_55 (.en(wire_305), .in(wire_8), .out(wire_83_18[15:0]));
  TC_Switch # (.UUID(64'd1287692551111612372 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_56 (.en(wire_110), .in(wire_421), .out(wire_83_19[15:0]));
  TC_Switch # (.UUID(64'd1141911395405296382 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_57 (.en(wire_218), .in({{8{1'b0}}, wire_199 }), .out(wire_83_20[15:0]));
  TC_Not # (.UUID(64'd3575339823787626444 ^ UUID), .BIT_WIDTH(64'd8)) Not8_58 (.in(wire_51[7:0]), .out(wire_199));
  TC_Rol # (.UUID(64'd2078177537373562034 ^ UUID), .BIT_WIDTH(64'd16)) Rol16_59 (.in(wire_51), .shift(wire_12[7:0]), .out(wire_421));
  TC_Shl # (.UUID(64'd4491813690601887022 ^ UUID), .BIT_WIDTH(64'd16)) Shl16_60 (.in(wire_51), .shift(wire_12[7:0]), .out(wire_76));
  TC_Shr # (.UUID(64'd4199576277751456538 ^ UUID), .BIT_WIDTH(64'd16)) Shr16_61 (.in(wire_51), .shift(wire_12[7:0]), .out(wire_353));
  TC_Xor # (.UUID(64'd1780129286836567965 ^ UUID), .BIT_WIDTH(64'd16)) Xor16_62 (.in0(wire_51), .in1(wire_12), .out(wire_106));
  TC_Or # (.UUID(64'd3629729579801707084 ^ UUID), .BIT_WIDTH(64'd16)) Or16_63 (.in0(wire_51), .in1(wire_12), .out(wire_288));
  TC_And # (.UUID(64'd3161317497787028707 ^ UUID), .BIT_WIDTH(64'd16)) And16_64 (.in0(wire_51), .in1(wire_12), .out(wire_390));
  TC_And # (.UUID(64'd381639147620396883 ^ UUID), .BIT_WIDTH(64'd8)) And8_65 (.in0(wire_272), .in1(wire_21[7:0]), .out(wire_235));
  TC_Or3 # (.UUID(64'd3488800466009071346 ^ UUID), .BIT_WIDTH(64'd1)) Or3_66 (.in0(wire_91), .in1(wire_88), .in2(wire_286), .out(wire_58));
  TC_Or # (.UUID(64'd800125638954551844 ^ UUID), .BIT_WIDTH(64'd1)) Or_67 (.in0(wire_221), .in1(wire_88), .out(wire_175));
  TC_Neg # (.UUID(64'd3923101654540497550 ^ UUID), .BIT_WIDTH(64'd16)) Neg16_68 (.in(wire_149), .out(wire_95));
  TC_Mux # (.UUID(64'd4466247896286800046 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_69 (.sel(wire_430), .in0(wire_95), .in1(wire_149), .out(wire_401));
  TC_Mux # (.UUID(64'd4573628848997923160 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_70 (.sel(wire_26), .in0({{8{1'b0}}, wire_437 }), .in1(wire_12), .out(wire_311));
  TC_Ashr # (.UUID(64'd2002805807653529301 ^ UUID), .BIT_WIDTH(64'd16)) Ashr16_71 (.in(wire_51), .shift(wire_12[7:0]), .out(wire_490));
  TC_Neg # (.UUID(64'd1410727121580829106 ^ UUID), .BIT_WIDTH(64'd16)) Neg16_72 (.in(wire_51), .out(wire_477));
  TC_Mul # (.UUID(64'd409697540344457906 ^ UUID), .BIT_WIDTH(64'd16)) DivMod16_73 (.in0(wire_51), .in1(wire_311), .out0(wire_289), .out1());
  TC_Mul # (.UUID(64'd4230356226461292418 ^ UUID), .BIT_WIDTH(64'd16)) Mul16_74 (.in0(wire_12), .in1(wire_51), .out0(wire_488), .out1());
  TC_Add # (.UUID(64'd1348307715225101930 ^ UUID), .BIT_WIDTH(64'd16)) Add16_75 (.in0(wire_401), .in1(wire_51), .ci(1'd0), .out(wire_348), .co());
  TC_Switch # (.UUID(64'd3604076901724081385 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_76 (.en(wire_192), .in(wire_477), .out(wire_83_9[15:0]));
  TC_Switch # (.UUID(64'd4522803089722429170 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_77 (.en(wire_26), .in(wire_289), .out(wire_83_11[15:0]));
  TC_Switch # (.UUID(64'd202434256468217393 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_78 (.en(wire_158), .in(wire_488), .out(wire_83_13[15:0]));
  TC_Switch # (.UUID(64'd981527730647914060 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_79 (.en(wire_58), .in(wire_348), .out(wire_83_15[15:0]));
  TC_IndexerByte # (.UUID(64'd4236276122307665751 ^ UUID), .INDEX(64'd0)) IndexerByte_80 (.in({{32{1'b0}}, wire_48 }), .out(wire_484));
  TC_Splitter8 # (.UUID(64'd4515369816812696921 ^ UUID)) Splitter8_81 (.in(wire_484), .out0(wire_286), .out1(wire_88), .out2(wire_158), .out3(wire_26), .out4(wire_192), .out5(wire_299), .out6(wire_221), .out7(wire_329));
  TC_Or # (.UUID(64'd3775589699623562439 ^ UUID), .BIT_WIDTH(64'd1)) Or_82 (.in0(wire_299), .in1(wire_221), .out(wire_91));
  TC_Or # (.UUID(64'd119900405875326486 ^ UUID), .BIT_WIDTH(64'd1)) Or_83 (.in0(wire_125), .in1(wire_228), .out(wire_183));
  TC_Add # (.UUID(64'd2771599484257026352 ^ UUID), .BIT_WIDTH(64'd16)) Add16_84 (.in0(wire_412), .in1(wire_303), .ci(1'd0), .out(wire_380), .co());
  TC_Mux # (.UUID(64'd1916750704823682311 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_85 (.sel(wire_72), .in0(wire_486), .in1(wire_155), .out(wire_217));
  TC_Switch # (.UUID(64'd110187611622282684 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_86 (.en(wire_43), .in(wire_233[15:0]), .out(wire_12_1));
  TC_Or # (.UUID(64'd1550338206798762433 ^ UUID), .BIT_WIDTH(64'd1)) Or_87 (.in0(wire_139), .in1(wire_141), .out(wire_137));
  TC_Switch # (.UUID(64'd1104805846581678264 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_88 (.en(wire_137), .in(wire_491[15:0]), .out(wire_51_0));
  TC_Or # (.UUID(64'd1973201053711173902 ^ UUID), .BIT_WIDTH(64'd1)) Or_89 (.in0(wire_141), .in1(wire_302), .out(wire_205));
  TC_And # (.UUID(64'd373051892767174731 ^ UUID), .BIT_WIDTH(64'd1)) And_90 (.in0(wire_265), .in1(wire_139), .out(wire_302));
  TC_Mux # (.UUID(64'd2189639269723513602 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_91 (.sel(wire_265), .in0(wire_173), .in1(wire_177), .out(wire_389));
  TC_Or3 # (.UUID(64'd4386189682368290849 ^ UUID), .BIT_WIDTH(64'd1)) Or3_92 (.in0(wire_141), .in1(wire_114), .in2(wire_265), .out(wire_284));
  TC_Nor # (.UUID(64'd3810192346818398090 ^ UUID), .BIT_WIDTH(64'd1)) Nor_93 (.in0(wire_284), .in1(wire_178), .out(wire_479));
  TC_Mux # (.UUID(64'd4107077995071586514 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_94 (.sel(wire_479), .in0(wire_389), .in1(wire_83[15:0]), .out(wire_56));
  TC_Switch # (.UUID(64'd1346494715147404059 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_95 (.en(wire_322), .in(wire_468), .out(wire_90_5));
  TC_Splitter8 # (.UUID(64'd3709071160935573773 ^ UUID)) Splitter8_96 (.in(wire_487), .out0(wire_229), .out1(wire_144), .out2(wire_145), .out3(wire_318), .out4(wire_413), .out5(wire_310), .out6(wire_322), .out7(wire_352));
  TC_Switch # (.UUID(64'd4272543595848591881 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_97 (.en(wire_144), .in(wire_478), .out(wire_90_4));
  TC_Switch # (.UUID(64'd2673250751246411725 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_98 (.en(wire_145), .in(wire_304), .out(wire_90_2));
  TC_Switch # (.UUID(64'd4158444071236719644 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_99 (.en(wire_318), .in(wire_258), .out(wire_90_0));
  TC_Switch # (.UUID(64'd1076960299062071464 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_100 (.en(wire_413), .in(wire_259), .out(wire_90_1));
  TC_Switch # (.UUID(64'd2871129963461955678 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_101 (.en(wire_310), .in(wire_449), .out(wire_90_3));
  TC_Switch # (.UUID(64'd1466219000736428262 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_102 (.en(wire_352), .in(wire_157), .out(wire_90_7));
  TC_LessU # (.UUID(64'd70784060852193480 ^ UUID), .BIT_WIDTH(64'd16)) LessU16_103 (.in0(wire_12), .in1(wire_51), .out(wire_157));
  TC_Or # (.UUID(64'd2633850717105506955 ^ UUID), .BIT_WIDTH(64'd1)) Or_104 (.in0(wire_157), .in1(wire_259), .out(wire_468));
  TC_Not # (.UUID(64'd2994142474806724920 ^ UUID), .BIT_WIDTH(64'd1)) Not_105 (.in(wire_259), .out(wire_449));
  TC_Equal # (.UUID(64'd4180772301230732474 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_106 (.in0(wire_51), .in1(wire_12), .out(wire_259));
  TC_LessU # (.UUID(64'd3216607671565821129 ^ UUID), .BIT_WIDTH(64'd16)) LessU16_107 (.in0(wire_51), .in1(wire_12), .out(wire_304));
  TC_Or # (.UUID(64'd1733367887190953979 ^ UUID), .BIT_WIDTH(64'd1)) Or_108 (.in0(wire_259), .in1(wire_304), .out(wire_258));
  TC_Equal # (.UUID(64'd2756161344151621510 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_109 (.in0({{8{1'b0}}, wire_425 }), .in1(wire_51), .out(wire_166));
  TC_Constant # (.UUID(64'd14059539423913175 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h0)) Constant8_110 (.out(wire_425));
  TC_Not # (.UUID(64'd2912282656104074477 ^ UUID), .BIT_WIDTH(64'd1)) Not_111 (.in(wire_166), .out(wire_478));
  TC_Switch # (.UUID(64'd338503895939097385 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_112 (.en(wire_229), .in(wire_166), .out(wire_90_6));
  TC_Switch # (.UUID(64'd2974250978505416008 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_113 (.en(wire_178), .in(wire_51), .out(wire_173));
  TC_Switch # (.UUID(64'd294942412853573551 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_114 (.en(wire_325), .in(wire_179), .out(wire_194_0));
  TC_Switch # (.UUID(64'd2530020128287448865 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_115 (.en(wire_241), .in(wire_123), .out(wire_194_1));
  TC_Not # (.UUID(64'd1944022449022311076 ^ UUID), .BIT_WIDTH(64'd1)) Not_116 (.in(wire_325), .out(wire_241));
  TC_Switch # (.UUID(64'd640117511591385720 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_117 (.en(wire_205), .in(wire_51), .out(wire_83_6[15:0]));
  TC_Clock # (.UUID(64'd473244454118914110 ^ UUID)) Clock_118 (.clk(clk), .rst(rst), .out(wire_325));
  TC_Switch # (.UUID(64'd3240978896697767469 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_119 (.en(wire_77), .in(wire_77), .out(wire_90_8));
  TC_Mux # (.UUID(64'd4327728578462997473 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_120 (.sel(wire_228), .in0(wire_217), .in1(wire_380), .out(wire_123));
  TC_Not # (.UUID(64'd2335834251709147674 ^ UUID), .BIT_WIDTH(64'd1)) Not_121 (.in(wire_138), .out(wire_295));
  TC_Switch # (.UUID(64'd1177966569030928993 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_122 (.en(wire_138), .in(wire_50), .out(wire_83_7[15:0]));
  TC_Switch # (.UUID(64'd4085565154656183842 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_123 (.en(wire_329), .in(wire_490), .out(wire_83_8[15:0]));
  TC_IndexerByte # (.UUID(64'd82359665637793120 ^ UUID), .INDEX(64'd2)) IndexerByte_124 (.in({{32{1'b0}}, wire_48 }), .out(wire_487));
  TC_Switch # (.UUID(64'd691486037870060392 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_125 (.en(wire_374), .in(wire_187), .out(wire_184));
  TC_IndexerBit # (.UUID(64'd1630189301439907508 ^ UUID), .INDEX(64'd4)) IndexerBit_126 (.in({{56{1'b0}}, wire_116 }), .out(wire_72));
  TC_IndexerBit # (.UUID(64'd2208263359456905046 ^ UUID), .INDEX(64'd5)) IndexerBit_127 (.in({{56{1'b0}}, wire_116 }), .out(wire_357));
  TC_IndexerByte # (.UUID(64'd2160584388702904456 ^ UUID), .INDEX(64'd3)) IndexerByte_128 (.in({{32{1'b0}}, wire_48 }), .out(wire_116));
  TC_Not # (.UUID(64'd904891828379418593 ^ UUID), .BIT_WIDTH(64'd1)) Not_129 (.in(wire_357), .out(wire_227));
  TC_Constant # (.UUID(64'd3538634162844758805 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hFF)) Constant8_130 (.out(wire_444));
  TC_Constant # (.UUID(64'd2648359173322761393 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hFE)) Constant8_131 (.out(wire_197));
  TC_Maker16 # (.UUID(64'd4168581648613032575 ^ UUID)) Maker16_132 (.in0(wire_444), .in1(wire_197), .out(wire_168));
  TC_Mux # (.UUID(64'd3090540701337537666 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_133 (.sel(wire_125), .in0(wire_366), .in1(wire_380), .out(wire_179));
  TC_Maker16 # (.UUID(64'd851087207377417069 ^ UUID)) Maker16_134 (.in0(wire_472), .in1(wire_239), .out(wire_303));
  TC_Constant # (.UUID(64'd381873739773538407 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hFF)) Constant8_135 (.out(wire_472));
  TC_Mux # (.UUID(64'd4592224200207251913 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_136 (.sel(wire_227), .in0(wire_207), .in1(wire_101), .out(wire_486));
  TC_Equal # (.UUID(64'd3099658865939077738 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_137 (.in0(wire_184), .in1(16'd0), .out(wire_215));
  TC_Not # (.UUID(64'd4471125710935676612 ^ UUID), .BIT_WIDTH(64'd1)) Not_138 (.in(wire_215), .out(wire_43));
  TC_IndexerBit # (.UUID(64'd460606693629125729 ^ UUID), .INDEX(64'd4)) IndexerBit_139 (.in({{56{1'b0}}, wire_103 }), .out(wire_265));
  TC_IndexerBit # (.UUID(64'd1499309531990315318 ^ UUID), .INDEX(64'd1)) IndexerBit_140 (.in({{56{1'b0}}, wire_103 }), .out(wire_114));
  TC_Or3 # (.UUID(64'd3834216222200410896 ^ UUID), .BIT_WIDTH(64'd1)) Or3_141 (.in0(wire_165), .in1(wire_485), .in2(wire_433), .out(wire_178));
  TC_IndexerBit # (.UUID(64'd345801079655292532 ^ UUID), .INDEX(64'd2)) IndexerBit_142 (.in({{56{1'b0}}, wire_103 }), .out(wire_485));
  TC_IndexerBit # (.UUID(64'd3857678701898454921 ^ UUID), .INDEX(64'd3)) IndexerBit_143 (.in({{56{1'b0}}, wire_103 }), .out(wire_165));
  TC_IndexerBit # (.UUID(64'd1094550749412879412 ^ UUID), .INDEX(64'd5)) IndexerBit_144 (.in({{56{1'b0}}, wire_103 }), .out(wire_141));
  TC_Not # (.UUID(64'd295801019876953925 ^ UUID), .BIT_WIDTH(64'd1)) Not_145 (.in(wire_481), .out(wire_146));
  TC_Equal # (.UUID(64'd3140328761418953014 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_146 (.in0(wire_179), .in1(16'd0), .out(wire_475));
  TC_Not # (.UUID(64'd4400946405007906585 ^ UUID), .BIT_WIDTH(64'd1)) Not_147 (.in(wire_266), .out(wire_139));
  TC_IndexerByte # (.UUID(64'd2633087214037843825 ^ UUID), .INDEX(64'd3)) IndexerByte_148 (.in({{32{1'b0}}, wire_48 }), .out(wire_103));
  TC_Equal # (.UUID(64'd2561182539117830921 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_149 (.in0(16'd0), .in1(wire_123), .out(wire_266));
  TC_IndexerBit # (.UUID(64'd2047893359182210890 ^ UUID), .INDEX(64'd0)) IndexerBit_150 (.in(wire_21), .out(wire_99));
  TC_IndexerBit # (.UUID(64'd3859884203355858265 ^ UUID), .INDEX(64'd1)) IndexerBit_151 (.in(wire_21), .out(wire_96));
  TC_IndexerBit # (.UUID(64'd4287739567158645737 ^ UUID), .INDEX(64'd2)) IndexerBit_152 (.in(wire_21), .out(wire_115));
  TC_IndexerBit # (.UUID(64'd777253982648504148 ^ UUID), .INDEX(64'd3)) IndexerBit_153 (.in(wire_21), .out(wire_296));
  TC_IndexerBit # (.UUID(64'd1771789865896455183 ^ UUID), .INDEX(64'd4)) IndexerBit_154 (.in(wire_21), .out(wire_5));
  TC_IndexerBit # (.UUID(64'd3105812192345802732 ^ UUID), .INDEX(64'd6)) IndexerBit_155 (.in(wire_21), .out(wire_307));
  TC_IndexerBit # (.UUID(64'd3077471030622112266 ^ UUID), .INDEX(64'd7)) IndexerBit_156 (.in(wire_21), .out(wire_373));
  TC_Not # (.UUID(64'd2159748274689718655 ^ UUID), .BIT_WIDTH(64'd1)) Not_157 (.in(wire_475), .out(wire_68));
  TC_Splitter16 # (.UUID(64'd1069070463351244943 ^ UUID)) Splitter16_158 (.in(wire_21[15:0]), .out0(), .out1(wire_385));
  TC_Switch # (.UUID(64'd3542778498052595836 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_159 (.en(wire_323), .in(wire_474[15:0]), .out(wire_83_2[15:0]));
  TC_Not # (.UUID(64'd944680686405816927 ^ UUID), .BIT_WIDTH(64'd1)) Not_160 (.in(wire_193), .out(wire_251));
  TC_Switch # (.UUID(64'd816465745217087424 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_161 (.en(wire_152), .in(wire_12), .out(wire_4));
  TC_Switch # (.UUID(64'd209623535459112064 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_162 (.en(wire_152), .in(wire_51), .out(wire_37));
  TC_And # (.UUID(64'd2522855677877010919 ^ UUID), .BIT_WIDTH(64'd1)) And_163 (.in0(wire_152), .in1(wire_410), .out(wire_323));
  TC_Equal # (.UUID(64'd2756262866884777429 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_164 (.in0(8'd0), .in1(wire_37[7:0]), .out(wire_410));
  TC_Equal # (.UUID(64'd1714264829042601315 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_165 (.in0(wire_385), .in1(wire_458), .out(wire_152));
  TC_Constant # (.UUID(64'd2907468583675662890 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_166 (.out(wire_458));
  TC_Mux # (.UUID(64'd2441497898305995710 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_167 (.sel(wire_72), .in0(wire_155), .in1(wire_207), .out(wire_366));
  TC_Switch # (.UUID(64'd3809517357945142409 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_168 (.en(wire_100), .in(wire_104[15:0]), .out(wire_25));
  TC_Not # (.UUID(64'd4003951151984714090 ^ UUID), .BIT_WIDTH(64'd1)) Not_169 (.in(wire_373), .out(wire_417));
  TC_IndexerBit # (.UUID(64'd1553590145675495351 ^ UUID), .INDEX(64'd5)) IndexerBit_170 (.in(wire_21), .out(wire_138));
  TC_Not # (.UUID(64'd3312304652180753239 ^ UUID), .BIT_WIDTH(64'd1)) Not_171 (.in(wire_307), .out(wire_374));
  TC_Constant # (.UUID(64'd2729531845625831067 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_172 (.out(wire_437));
  TC_Not # (.UUID(64'd2538698523318428916 ^ UUID), .BIT_WIDTH(64'd1)) Not_173 (.in(wire_175), .out(wire_430));
  TC_Constant # (.UUID(64'd2179489257373318160 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_174 (.out(wire_273));
  TC_Mux # (.UUID(64'd2429066787419951843 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_175 (.sel(wire_91), .in0(wire_12), .in1({{8{1'b0}}, wire_273 }), .out(wire_149));
  TC_Switch # (.UUID(64'd391371808230282023 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_176 (.en(wire_203), .in(wire_195), .out(wire_267));
  TC_Constant # (.UUID(64'd2691125905525222303 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1F)) Constant8_177 (.out(wire_272));
  TC_IndexerByte # (.UUID(64'd2112170900386343144 ^ UUID), .INDEX(64'd3)) IndexerByte_178 (.in({{32{1'b0}}, wire_48 }), .out(wire_164));
  TC_IndexerBit # (.UUID(64'd2727080739164391000 ^ UUID), .INDEX(64'd6)) IndexerBit_179 (.in({{56{1'b0}}, wire_164 }), .out(wire_301));
  TC_Switch # (.UUID(64'd2160087561000370162 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_180 (.en(wire_301), .in(wire_301), .out(wire_90_9));
  TC_Switch # (.UUID(64'd592302940647155691 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_181 (.en(wire_426), .in({{15{1'b0}}, wire_394 }), .out(wire_83_5[15:0]));
  TC_Or # (.UUID(64'd3278179513885088927 ^ UUID), .BIT_WIDTH(64'd1)) Or_182 (.in0(wire_426), .in1(wire_387), .out(wire_334));
  TC_Equal # (.UUID(64'd4033274235037801114 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_183 (.in0(wire_467), .in1(wire_245), .out(wire_426));
  TC_Not # (.UUID(64'd1697593568395826930 ^ UUID), .BIT_WIDTH(64'd1)) Not_184 (.in(wire_387), .out(wire_386));
  TC_Splitter16 # (.UUID(64'd962308306064647197 ^ UUID)) Splitter16_185 (.in(wire_21[15:0]), .out0(), .out1(wire_467));
  TC_Constant # (.UUID(64'd3037869375563223000 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h2)) Constant8_186 (.out(wire_245));
  TC_DelayLine # (.UUID(64'd4275385609773382257 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_187 (.clk(clk), .rst(rst), .in(wire_291), .out(wire_387));
  TC_Switch # (.UUID(64'd1286392688347840013 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_188 (.en(wire_386), .in(wire_334), .out(wire_291));
  TC_Splitter16 # (.UUID(64'd815166994044352782 ^ UUID)) Splitter16_189 (.in(wire_21[15:0]), .out0(), .out1(wire_202));
  TC_IndexerByte # (.UUID(64'd4056757385308142069 ^ UUID), .INDEX(64'd1)) IndexerByte_190 (.in(wire_359), .out(wire_471));
  TC_IndexerByte # (.UUID(64'd4445007758314830950 ^ UUID), .INDEX(64'd0)) IndexerByte_191 (.in(wire_359), .out(wire_253));
  TC_Maker16 # (.UUID(64'd1879612468053834457 ^ UUID)) Maker16_192 (.in0(wire_253), .in1(wire_471), .out(wire_395));
  TC_Switch # (.UUID(64'd220823607166135876 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_193 (.en(wire_94), .in(wire_395), .out(wire_83_0[15:0]));
  TC_Equal # (.UUID(64'd3724760983101447498 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_194 (.in0(wire_202), .in1(wire_416), .out(wire_94));
  TC_Constant # (.UUID(64'd1337227511337026411 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h3)) Constant8_195 (.out(wire_416));
  TC_Timing # (.UUID(64'd2799049267103079424 ^ UUID)) Timing_196 (.en(wire_94), .out(wire_359));
  TC_Program # (.UUID(64'd3721980137216604240 ^ UUID), .WORD_WIDTH(64'd8), .DEFAULT_FILE_NAME("Program_33A7213703DAF850.w8.bin"), .ARG_SIG("Program_33A7213703DAF850=%s")) Program_197 (.clk(clk), .rst(rst), .address(wire_51), .out0(wire_294), .out1(), .out2(), .out3());
  TC_Splitter16 # (.UUID(64'd4461787469973933422 ^ UUID)) Splitter16_198 (.in(wire_21[15:0]), .out0(), .out1(wire_476));
  TC_Equal # (.UUID(64'd1988770091565985332 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_199 (.in0(wire_476), .in1(wire_35), .out(wire_181));
  TC_Constant # (.UUID(64'd2565543928344869306 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h5)) Constant8_200 (.out(wire_35));
  TC_Switch # (.UUID(64'd4105771623231641306 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_201 (.en(wire_181), .in(wire_294[15:0]), .out(wire_83_4[15:0]));
  TC_Equal # (.UUID(64'd551722571517782638 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_202 (.in0(16'd0), .in1(wire_37), .out(wire_193));
  TC_Register # (.UUID(64'd4364107987795409853 ^ UUID), .BIT_WIDTH(64'd16)) Register16_203 (.clk(clk), .rst(rst), .load(wire_183), .save(wire_183), .in(wire_312), .out(wire_74));
  TC_Constant # (.UUID(64'd1415884859697557611 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_204 (.out(wire_108));
  TC_IndexerBit # (.UUID(64'd535377880148297947 ^ UUID), .INDEX(64'd3)) IndexerBit_205 (.in({{56{1'b0}}, wire_116 }), .out(wire_228));
  TC_Register # (.UUID(64'd2160598746671012754 ^ UUID), .BIT_WIDTH(64'd16)) Register16_206 (.clk(clk), .rst(rst), .load(wire_77), .save(wire_77), .in(wire_136), .out(wire_206));
  TC_Add # (.UUID(64'd1442806402229030427 ^ UUID), .BIT_WIDTH(64'd16)) Add16_207 (.in0(wire_298), .in1(wire_168), .ci(1'd0), .out(wire_207), .co());
  TC_Or # (.UUID(64'd2188959817660993009 ^ UUID), .BIT_WIDTH(64'd1)) Or_208 (.in0(wire_72), .in1(wire_357), .out(wire_77));
  TC_IndexerBit # (.UUID(64'd3588176080026118662 ^ UUID), .INDEX(64'd2)) IndexerBit_209 (.in({{56{1'b0}}, wire_116 }), .out(wire_125));
  TC_Mux # (.UUID(64'd4063471477342436371 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_210 (.sel(wire_357), .in0(wire_346), .in1(wire_206), .out(wire_298));
  TC_Mux # (.UUID(64'd527759690959107192 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_211 (.sel(wire_228), .in0(wire_392), .in1(wire_74), .out(wire_412));
  TC_Switch # (.UUID(64'd1362725833065582892 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_212 (.en(wire_125), .in(wire_312), .out(wire_392));
  TC_Switch # (.UUID(64'd1756831740426205013 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_213 (.en(wire_72), .in(wire_136), .out(wire_346));
  TC_Add # (.UUID(64'd2930665708224337659 ^ UUID), .BIT_WIDTH(64'd16)) Add16_214 (.in0(wire_74), .in1(wire_293), .ci(1'd0), .out(wire_312), .co());
  TC_Constant # (.UUID(64'd3137150186803814383 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hF0)) Constant8_215 (.out(wire_239));
  TC_Add # (.UUID(64'd432537638553101254 ^ UUID), .BIT_WIDTH(64'd16)) Add16_216 (.in0(wire_206), .in1(wire_190), .ci(1'd0), .out(wire_136), .co());
  TC_IndexerBit # (.UUID(64'd561707948535025464 ^ UUID), .INDEX(64'd4)) IndexerBit_217 (.in({{56{1'b0}}, wire_116 }), .out(wire_268));
  TC_Constant # (.UUID(64'd1695694096694981758 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_218 (.out(wire_344));
  TC_IndexerBit # (.UUID(64'd2331812482237933900 ^ UUID), .INDEX(64'd0)) IndexerBit_219 (.in({{56{1'b0}}, wire_269 }), .out(wire_433));
  TC_Neg # (.UUID(64'd1821476619534246961 ^ UUID), .BIT_WIDTH(64'd16)) Neg16_220 (.in({{8{1'b0}}, wire_344 }), .out(wire_439));
  TC_Mux # (.UUID(64'd1539425850473868597 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_221 (.sel(wire_268), .in0(wire_439), .in1({{8{1'b0}}, wire_344 }), .out(wire_190));
  TC_Mux # (.UUID(64'd3572805427243657698 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_222 (.sel(wire_125), .in0(wire_80), .in1({{8{1'b0}}, wire_108 }), .out(wire_293));
  TC_Neg # (.UUID(64'd2090057048615449572 ^ UUID), .BIT_WIDTH(64'd16)) Neg16_223 (.in({{8{1'b0}}, wire_108 }), .out(wire_80));
  TC_IOSwitch # (.UUID(64'd2846053541171193881 ^ UUID), .BIT_WIDTH(64'd8)) LevelOutputArch_224 (.in(wire_51[7:0]), .en(wire_338), .out(arch_output_value));
  TC_Switch # (.UUID(64'd210661621448949326 ^ UUID), .BIT_WIDTH(64'd8)) LevelInputArch_225 (.en(wire_398), .in(arch_input_value), .out(wire_83_3[7:0]));
  TC_Splitter16 # (.UUID(64'd2775342692045340835 ^ UUID)) Splitter16_226 (.in(wire_21[15:0]), .out0(), .out1(wire_320));
  TC_Equal # (.UUID(64'd4532639728004948159 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_227 (.in0(wire_320), .in1(wire_214), .out(wire_261));
  TC_Equal # (.UUID(64'd3745587913460272427 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_228 (.in0(wire_419), .in1(wire_320), .out(wire_400));
  TC_Constant # (.UUID(64'd951998662890801082 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6)) Constant8_229 (.out(wire_419));
  TC_Constant # (.UUID(64'd2262634952183580731 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7)) Constant8_230 (.out(wire_214));
  TC_Switch # (.UUID(64'd1419008802292368204 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_231 (.en(wire_237), .in(wire_400), .out(wire_398));
  TC_Clock # (.UUID(64'd150335021447124340 ^ UUID)) Clock_232 (.clk(clk), .rst(rst), .out(wire_237));
  TC_Switch # (.UUID(64'd3781955660154943019 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_233 (.en(wire_415), .in(wire_261), .out(wire_338));
  TC_Not # (.UUID(64'd248590985388437467 ^ UUID), .BIT_WIDTH(64'd1)) Not_234 (.in(wire_237), .out(wire_415));
  TC_RamDualLoad # (.UUID(64'd1162091816344660036 ^ UUID), .WORD_WIDTH(64'd16), .WORD_COUNT(64'd65536)) RamDualLoad_235 (.clk(clk), .rst(rst), .load0(wire_139), .save(wire_68), .address0({{16{1'b0}}, wire_194 }), .in({{48{1'b0}}, wire_56 }), .load1(wire_43), .address1({{16{1'b0}}, wire_184 }), .out0(wire_491), .out1(wire_233));
  TC_Ram # (.UUID(64'd2071862132571227302 ^ UUID), .WORD_WIDTH(64'd16), .WORD_COUNT(64'd65536)) Ram_236 (.clk(clk), .rst(rst), .load(wire_193), .save(wire_251), .address({{16{1'b0}}, wire_4 }), .in0({{48{1'b0}}, wire_37 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_474), .out1(), .out2(), .out3());
  TC_FileLoader # (.UUID(64'd1149854990232492044 ^ UUID), .DEFAULT_FILE_NAME("image.dat")) FileLoader_237 (.clk(clk), .rst(rst), .en(wire_264), .address({{48{1'b0}}, wire_51 }), .out(wire_83_1));
  TC_Splitter16 # (.UUID(64'd2684349980131024015 ^ UUID)) Splitter16_238 (.in(wire_21[15:0]), .out0(), .out1(wire_431));
  TC_Equal # (.UUID(64'd4369488988257915881 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_239 (.in0(wire_431), .in1(wire_436), .out(wire_264));
  TC_Constant # (.UUID(64'd3823619217162964047 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hA)) Constant8_240 (.out(wire_436));
  TC_Ror # (.UUID(64'd445352019034615982 ^ UUID), .BIT_WIDTH(64'd16)) Ror16_241 (.in(wire_51), .shift(wire_12[7:0]), .out(wire_8));
  TC_DotMatrixDisplay # (.UUID(64'd194337641353170009 ^ UUID)) DotMatrixDisplay_242 (.clk(clk), .rst(rst), .en_y(wire_111[0:0]), .en_x(wire_38[0:0]), .color_info(wire_111), .pixel_info(wire_38));
  TC_DotMatrixDisplay # (.UUID(64'd2571677606765972402 ^ UUID)) DotMatrixDisplay_243 (.clk(clk), .rst(rst), .en_y(wire_6[0:0]), .en_x(wire_38[0:0]), .color_info(wire_6), .pixel_info(wire_38));
  TC_DotMatrixDisplay # (.UUID(64'd138839058832846553 ^ UUID)) DotMatrixDisplay_244 (.clk(clk), .rst(rst), .en_y(wire_67[0:0]), .en_x(wire_38[0:0]), .color_info(wire_67), .pixel_info(wire_38));
  TC_DotMatrixDisplay # (.UUID(64'd3101733260034986425 ^ UUID)) DotMatrixDisplay_245 (.clk(clk), .rst(rst), .en_y(wire_44[0:0]), .en_x(wire_38[0:0]), .color_info(wire_44), .pixel_info(wire_38));
  TC_DotMatrixDisplay # (.UUID(64'd4009925455146135119 ^ UUID)) DotMatrixDisplay_246 (.clk(clk), .rst(rst), .en_y(wire_49[0:0]), .en_x(wire_38[0:0]), .color_info(wire_49), .pixel_info(wire_38));
  TC_DotMatrixDisplay # (.UUID(64'd4277063417422545180 ^ UUID)) DotMatrixDisplay_247 (.clk(clk), .rst(rst), .en_y(wire_71[0:0]), .en_x(wire_38[0:0]), .color_info(wire_71), .pixel_info(wire_38));
  TC_DotMatrixDisplay # (.UUID(64'd58773507439597400 ^ UUID)) DotMatrixDisplay_248 (.clk(clk), .rst(rst), .en_y(wire_1[0:0]), .en_x(wire_38[0:0]), .color_info(wire_1), .pixel_info(wire_38));
  TC_DotMatrixDisplay # (.UUID(64'd3718278364047458166 ^ UUID)) DotMatrixDisplay_249 (.clk(clk), .rst(rst), .en_y(wire_111[0:0]), .en_x(wire_46[0:0]), .color_info(wire_111), .pixel_info(wire_46));
  TC_DotMatrixDisplay # (.UUID(64'd3828063013731251984 ^ UUID)) DotMatrixDisplay_250 (.clk(clk), .rst(rst), .en_y(wire_6[0:0]), .en_x(wire_46[0:0]), .color_info(wire_6), .pixel_info(wire_46));
  TC_DotMatrixDisplay # (.UUID(64'd3173625762873083734 ^ UUID)) DotMatrixDisplay_251 (.clk(clk), .rst(rst), .en_y(wire_67[0:0]), .en_x(wire_46[0:0]), .color_info(wire_67), .pixel_info(wire_46));
  TC_DotMatrixDisplay # (.UUID(64'd4159247278947979257 ^ UUID)) DotMatrixDisplay_252 (.clk(clk), .rst(rst), .en_y(wire_44[0:0]), .en_x(wire_46[0:0]), .color_info(wire_44), .pixel_info(wire_46));
  TC_DotMatrixDisplay # (.UUID(64'd841450751213016891 ^ UUID)) DotMatrixDisplay_253 (.clk(clk), .rst(rst), .en_y(wire_49[0:0]), .en_x(wire_46[0:0]), .color_info(wire_49), .pixel_info(wire_46));
  TC_DotMatrixDisplay # (.UUID(64'd18461418125437468 ^ UUID)) DotMatrixDisplay_254 (.clk(clk), .rst(rst), .en_y(wire_71[0:0]), .en_x(wire_46[0:0]), .color_info(wire_71), .pixel_info(wire_46));
  TC_DotMatrixDisplay # (.UUID(64'd1499808489686266316 ^ UUID)) DotMatrixDisplay_255 (.clk(clk), .rst(rst), .en_y(wire_1[0:0]), .en_x(wire_46[0:0]), .color_info(wire_1), .pixel_info(wire_46));
  TC_DotMatrixDisplay # (.UUID(64'd1491673485310828437 ^ UUID)) DotMatrixDisplay_256 (.clk(clk), .rst(rst), .en_y(wire_111[0:0]), .en_x(wire_16[0:0]), .color_info(wire_111), .pixel_info(wire_16));
  TC_DotMatrixDisplay # (.UUID(64'd3056379081757526387 ^ UUID)) DotMatrixDisplay_257 (.clk(clk), .rst(rst), .en_y(wire_6[0:0]), .en_x(wire_16[0:0]), .color_info(wire_6), .pixel_info(wire_16));
  TC_DotMatrixDisplay # (.UUID(64'd937174553272161025 ^ UUID)) DotMatrixDisplay_258 (.clk(clk), .rst(rst), .en_y(wire_67[0:0]), .en_x(wire_16[0:0]), .color_info(wire_67), .pixel_info(wire_16));
  TC_DotMatrixDisplay # (.UUID(64'd3051308917649846056 ^ UUID)) DotMatrixDisplay_259 (.clk(clk), .rst(rst), .en_y(wire_44[0:0]), .en_x(wire_16[0:0]), .color_info(wire_44), .pixel_info(wire_16));
  TC_DotMatrixDisplay # (.UUID(64'd2751084514686000524 ^ UUID)) DotMatrixDisplay_260 (.clk(clk), .rst(rst), .en_y(wire_49[0:0]), .en_x(wire_16[0:0]), .color_info(wire_49), .pixel_info(wire_16));
  TC_DotMatrixDisplay # (.UUID(64'd1256511526243769959 ^ UUID)) DotMatrixDisplay_261 (.clk(clk), .rst(rst), .en_y(wire_71[0:0]), .en_x(wire_16[0:0]), .color_info(wire_71), .pixel_info(wire_16));
  TC_DotMatrixDisplay # (.UUID(64'd2075225446636166702 ^ UUID)) DotMatrixDisplay_262 (.clk(clk), .rst(rst), .en_y(wire_1[0:0]), .en_x(wire_16[0:0]), .color_info(wire_1), .pixel_info(wire_16));
  TC_DotMatrixDisplay # (.UUID(64'd2738388019733878846 ^ UUID)) DotMatrixDisplay_263 (.clk(clk), .rst(rst), .en_y(wire_111[0:0]), .en_x(wire_11[0:0]), .color_info(wire_111), .pixel_info(wire_11));
  TC_DotMatrixDisplay # (.UUID(64'd1346613707047915800 ^ UUID)) DotMatrixDisplay_264 (.clk(clk), .rst(rst), .en_y(wire_6[0:0]), .en_x(wire_11[0:0]), .color_info(wire_6), .pixel_info(wire_11));
  TC_DotMatrixDisplay # (.UUID(64'd4578970333081576098 ^ UUID)) DotMatrixDisplay_265 (.clk(clk), .rst(rst), .en_y(wire_67[0:0]), .en_x(wire_11[0:0]), .color_info(wire_67), .pixel_info(wire_11));
  TC_DotMatrixDisplay # (.UUID(64'd2397741494846183167 ^ UUID)) DotMatrixDisplay_266 (.clk(clk), .rst(rst), .en_y(wire_44[0:0]), .en_x(wire_11[0:0]), .color_info(wire_44), .pixel_info(wire_11));
  TC_DotMatrixDisplay # (.UUID(64'd2638784560376988785 ^ UUID)) DotMatrixDisplay_267 (.clk(clk), .rst(rst), .en_y(wire_49[0:0]), .en_x(wire_11[0:0]), .color_info(wire_49), .pixel_info(wire_11));
  TC_DotMatrixDisplay # (.UUID(64'd4528084328396190170 ^ UUID)) DotMatrixDisplay_268 (.clk(clk), .rst(rst), .en_y(wire_71[0:0]), .en_x(wire_11[0:0]), .color_info(wire_71), .pixel_info(wire_11));
  TC_DotMatrixDisplay # (.UUID(64'd3851842690265338608 ^ UUID)) DotMatrixDisplay_269 (.clk(clk), .rst(rst), .en_y(wire_1[0:0]), .en_x(wire_11[0:0]), .color_info(wire_1), .pixel_info(wire_11));
  TC_DotMatrixDisplay # (.UUID(64'd4007736008231897574 ^ UUID)) DotMatrixDisplay_270 (.clk(clk), .rst(rst), .en_y(wire_111[0:0]), .en_x(wire_65[0:0]), .color_info(wire_111), .pixel_info(wire_65));
  TC_DotMatrixDisplay # (.UUID(64'd3826021121295671528 ^ UUID)) DotMatrixDisplay_271 (.clk(clk), .rst(rst), .en_y(wire_6[0:0]), .en_x(wire_65[0:0]), .color_info(wire_6), .pixel_info(wire_65));
  TC_DotMatrixDisplay # (.UUID(64'd4588979816491789595 ^ UUID)) DotMatrixDisplay_272 (.clk(clk), .rst(rst), .en_y(wire_67[0:0]), .en_x(wire_65[0:0]), .color_info(wire_67), .pixel_info(wire_65));
  TC_DotMatrixDisplay # (.UUID(64'd471994117323042265 ^ UUID)) DotMatrixDisplay_273 (.clk(clk), .rst(rst), .en_y(wire_44[0:0]), .en_x(wire_65[0:0]), .color_info(wire_44), .pixel_info(wire_65));
  TC_DotMatrixDisplay # (.UUID(64'd3038285795447948478 ^ UUID)) DotMatrixDisplay_274 (.clk(clk), .rst(rst), .en_y(wire_49[0:0]), .en_x(wire_65[0:0]), .color_info(wire_49), .pixel_info(wire_65));
  TC_DotMatrixDisplay # (.UUID(64'd4581525392239126243 ^ UUID)) DotMatrixDisplay_275 (.clk(clk), .rst(rst), .en_y(wire_71[0:0]), .en_x(wire_65[0:0]), .color_info(wire_71), .pixel_info(wire_65));
  TC_DotMatrixDisplay # (.UUID(64'd1436097369683470840 ^ UUID)) DotMatrixDisplay_276 (.clk(clk), .rst(rst), .en_y(wire_1[0:0]), .en_x(wire_65[0:0]), .color_info(wire_1), .pixel_info(wire_65));
  TC_DotMatrixDisplay # (.UUID(64'd499728826686780779 ^ UUID)) DotMatrixDisplay_277 (.clk(clk), .rst(rst), .en_y(wire_111[0:0]), .en_x(wire_7[0:0]), .color_info(wire_111), .pixel_info(wire_7));
  TC_DotMatrixDisplay # (.UUID(64'd1543247313219277311 ^ UUID)) DotMatrixDisplay_278 (.clk(clk), .rst(rst), .en_y(wire_6[0:0]), .en_x(wire_7[0:0]), .color_info(wire_6), .pixel_info(wire_7));
  TC_DotMatrixDisplay # (.UUID(64'd1693499669572890407 ^ UUID)) DotMatrixDisplay_279 (.clk(clk), .rst(rst), .en_y(wire_67[0:0]), .en_x(wire_7[0:0]), .color_info(wire_67), .pixel_info(wire_7));
  TC_DotMatrixDisplay # (.UUID(64'd647796916272613197 ^ UUID)) DotMatrixDisplay_280 (.clk(clk), .rst(rst), .en_y(wire_44[0:0]), .en_x(wire_7[0:0]), .color_info(wire_44), .pixel_info(wire_7));
  TC_DotMatrixDisplay # (.UUID(64'd2848040708874525941 ^ UUID)) DotMatrixDisplay_281 (.clk(clk), .rst(rst), .en_y(wire_49[0:0]), .en_x(wire_7[0:0]), .color_info(wire_49), .pixel_info(wire_7));
  TC_DotMatrixDisplay # (.UUID(64'd3459540269725230160 ^ UUID)) DotMatrixDisplay_282 (.clk(clk), .rst(rst), .en_y(wire_71[0:0]), .en_x(wire_7[0:0]), .color_info(wire_71), .pixel_info(wire_7));
  TC_DotMatrixDisplay # (.UUID(64'd3827924278582584392 ^ UUID)) DotMatrixDisplay_283 (.clk(clk), .rst(rst), .en_y(wire_1[0:0]), .en_x(wire_7[0:0]), .color_info(wire_1), .pixel_info(wire_7));
  TC_DotMatrixDisplay # (.UUID(64'd3058896873561121055 ^ UUID)) DotMatrixDisplay_284 (.clk(clk), .rst(rst), .en_y(wire_111[0:0]), .en_x(wire_52[0:0]), .color_info(wire_111), .pixel_info(wire_52));
  TC_DotMatrixDisplay # (.UUID(64'd640281640035612674 ^ UUID)) DotMatrixDisplay_285 (.clk(clk), .rst(rst), .en_y(wire_6[0:0]), .en_x(wire_52[0:0]), .color_info(wire_6), .pixel_info(wire_52));
  TC_DotMatrixDisplay # (.UUID(64'd53313000373404008 ^ UUID)) DotMatrixDisplay_286 (.clk(clk), .rst(rst), .en_y(wire_67[0:0]), .en_x(wire_52[0:0]), .color_info(wire_67), .pixel_info(wire_52));
  TC_DotMatrixDisplay # (.UUID(64'd1293625241450709160 ^ UUID)) DotMatrixDisplay_287 (.clk(clk), .rst(rst), .en_y(wire_44[0:0]), .en_x(wire_52[0:0]), .color_info(wire_44), .pixel_info(wire_52));
  TC_DotMatrixDisplay # (.UUID(64'd1548081783831727021 ^ UUID)) DotMatrixDisplay_288 (.clk(clk), .rst(rst), .en_y(wire_49[0:0]), .en_x(wire_52[0:0]), .color_info(wire_49), .pixel_info(wire_52));
  TC_DotMatrixDisplay # (.UUID(64'd1196844806900845054 ^ UUID)) DotMatrixDisplay_289 (.clk(clk), .rst(rst), .en_y(wire_71[0:0]), .en_x(wire_52[0:0]), .color_info(wire_71), .pixel_info(wire_52));
  TC_DotMatrixDisplay # (.UUID(64'd304219024799832638 ^ UUID)) DotMatrixDisplay_290 (.clk(clk), .rst(rst), .en_y(wire_1[0:0]), .en_x(wire_52[0:0]), .color_info(wire_1), .pixel_info(wire_52));
  TC_DotMatrixDisplay # (.UUID(64'd3495013800602512637 ^ UUID)) DotMatrixDisplay_291 (.clk(clk), .rst(rst), .en_y(wire_111[0:0]), .en_x(wire_41[0:0]), .color_info(wire_111), .pixel_info(wire_41));
  TC_DotMatrixDisplay # (.UUID(64'd1115162128073258755 ^ UUID)) DotMatrixDisplay_292 (.clk(clk), .rst(rst), .en_y(wire_6[0:0]), .en_x(wire_41[0:0]), .color_info(wire_6), .pixel_info(wire_41));
  TC_DotMatrixDisplay # (.UUID(64'd4145032985905828907 ^ UUID)) DotMatrixDisplay_293 (.clk(clk), .rst(rst), .en_y(wire_67[0:0]), .en_x(wire_41[0:0]), .color_info(wire_67), .pixel_info(wire_41));
  TC_DotMatrixDisplay # (.UUID(64'd3507470446193958289 ^ UUID)) DotMatrixDisplay_294 (.clk(clk), .rst(rst), .en_y(wire_44[0:0]), .en_x(wire_41[0:0]), .color_info(wire_44), .pixel_info(wire_41));
  TC_DotMatrixDisplay # (.UUID(64'd1946383192464286856 ^ UUID)) DotMatrixDisplay_295 (.clk(clk), .rst(rst), .en_y(wire_49[0:0]), .en_x(wire_41[0:0]), .color_info(wire_49), .pixel_info(wire_41));
  TC_DotMatrixDisplay # (.UUID(64'd3575583628724029497 ^ UUID)) DotMatrixDisplay_296 (.clk(clk), .rst(rst), .en_y(wire_71[0:0]), .en_x(wire_41[0:0]), .color_info(wire_71), .pixel_info(wire_41));
  TC_DotMatrixDisplay # (.UUID(64'd1888768381846068356 ^ UUID)) DotMatrixDisplay_297 (.clk(clk), .rst(rst), .en_y(wire_1[0:0]), .en_x(wire_41[0:0]), .color_info(wire_1), .pixel_info(wire_41));
  TC_DotMatrixDisplay # (.UUID(64'd21752811922838239 ^ UUID)) DotMatrixDisplay_298 (.clk(clk), .rst(rst), .en_y(wire_111[0:0]), .en_x(wire_59[0:0]), .color_info(wire_111), .pixel_info(wire_59));
  TC_DotMatrixDisplay # (.UUID(64'd4252941668864125794 ^ UUID)) DotMatrixDisplay_299 (.clk(clk), .rst(rst), .en_y(wire_6[0:0]), .en_x(wire_59[0:0]), .color_info(wire_6), .pixel_info(wire_59));
  TC_DotMatrixDisplay # (.UUID(64'd2630952713397965447 ^ UUID)) DotMatrixDisplay_300 (.clk(clk), .rst(rst), .en_y(wire_67[0:0]), .en_x(wire_59[0:0]), .color_info(wire_67), .pixel_info(wire_59));
  TC_DotMatrixDisplay # (.UUID(64'd1603899630562403024 ^ UUID)) DotMatrixDisplay_301 (.clk(clk), .rst(rst), .en_y(wire_44[0:0]), .en_x(wire_59[0:0]), .color_info(wire_44), .pixel_info(wire_59));
  TC_DotMatrixDisplay # (.UUID(64'd2334824276736164064 ^ UUID)) DotMatrixDisplay_302 (.clk(clk), .rst(rst), .en_y(wire_49[0:0]), .en_x(wire_59[0:0]), .color_info(wire_49), .pixel_info(wire_59));
  TC_DotMatrixDisplay # (.UUID(64'd1944255304492587035 ^ UUID)) DotMatrixDisplay_303 (.clk(clk), .rst(rst), .en_y(wire_71[0:0]), .en_x(wire_59[0:0]), .color_info(wire_71), .pixel_info(wire_59));
  TC_DotMatrixDisplay # (.UUID(64'd3651443781059433220 ^ UUID)) DotMatrixDisplay_304 (.clk(clk), .rst(rst), .en_y(wire_1[0:0]), .en_x(wire_59[0:0]), .color_info(wire_1), .pixel_info(wire_59));
  TC_DotMatrixDisplay # (.UUID(64'd1676036236038663672 ^ UUID)) DotMatrixDisplay_305 (.clk(clk), .rst(rst), .en_y(wire_111[0:0]), .en_x(wire_30[0:0]), .color_info(wire_111), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd4189338739261535131 ^ UUID)) DotMatrixDisplay_306 (.clk(clk), .rst(rst), .en_y(wire_6[0:0]), .en_x(wire_30[0:0]), .color_info(wire_6), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd1091606415562326239 ^ UUID)) DotMatrixDisplay_307 (.clk(clk), .rst(rst), .en_y(wire_67[0:0]), .en_x(wire_30[0:0]), .color_info(wire_67), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd3980583843893868044 ^ UUID)) DotMatrixDisplay_308 (.clk(clk), .rst(rst), .en_y(wire_44[0:0]), .en_x(wire_30[0:0]), .color_info(wire_44), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd2842701554999032512 ^ UUID)) DotMatrixDisplay_309 (.clk(clk), .rst(rst), .en_y(wire_49[0:0]), .en_x(wire_30[0:0]), .color_info(wire_49), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd674998757530414630 ^ UUID)) DotMatrixDisplay_310 (.clk(clk), .rst(rst), .en_y(wire_71[0:0]), .en_x(wire_30[0:0]), .color_info(wire_71), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd1659403064194610874 ^ UUID)) DotMatrixDisplay_311 (.clk(clk), .rst(rst), .en_y(wire_1[0:0]), .en_x(wire_30[0:0]), .color_info(wire_1), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd2385476680905484428 ^ UUID)) DotMatrixDisplay_312 (.clk(clk), .rst(rst), .en_y(wire_111[0:0]), .en_x(wire_57[0:0]), .color_info(wire_111), .pixel_info(wire_57));
  TC_DotMatrixDisplay # (.UUID(64'd1405081695436727065 ^ UUID)) DotMatrixDisplay_313 (.clk(clk), .rst(rst), .en_y(wire_6[0:0]), .en_x(wire_57[0:0]), .color_info(wire_6), .pixel_info(wire_57));
  TC_DotMatrixDisplay # (.UUID(64'd996918915708390693 ^ UUID)) DotMatrixDisplay_314 (.clk(clk), .rst(rst), .en_y(wire_67[0:0]), .en_x(wire_57[0:0]), .color_info(wire_67), .pixel_info(wire_57));
  TC_DotMatrixDisplay # (.UUID(64'd2606453016393261708 ^ UUID)) DotMatrixDisplay_315 (.clk(clk), .rst(rst), .en_y(wire_44[0:0]), .en_x(wire_57[0:0]), .color_info(wire_44), .pixel_info(wire_57));
  TC_DotMatrixDisplay # (.UUID(64'd128040519194868715 ^ UUID)) DotMatrixDisplay_316 (.clk(clk), .rst(rst), .en_y(wire_49[0:0]), .en_x(wire_57[0:0]), .color_info(wire_49), .pixel_info(wire_57));
  TC_DotMatrixDisplay # (.UUID(64'd4546969349354631509 ^ UUID)) DotMatrixDisplay_317 (.clk(clk), .rst(rst), .en_y(wire_71[0:0]), .en_x(wire_57[0:0]), .color_info(wire_71), .pixel_info(wire_57));
  TC_DotMatrixDisplay # (.UUID(64'd1811149671421223324 ^ UUID)) DotMatrixDisplay_318 (.clk(clk), .rst(rst), .en_y(wire_1[0:0]), .en_x(wire_57[0:0]), .color_info(wire_1), .pixel_info(wire_57));
  TC_DotMatrixDisplay # (.UUID(64'd526846705743514459 ^ UUID)) DotMatrixDisplay_319 (.clk(clk), .rst(rst), .en_y(wire_111[0:0]), .en_x(wire_33[0:0]), .color_info(wire_111), .pixel_info(wire_33));
  TC_DotMatrixDisplay # (.UUID(64'd2410506663546344078 ^ UUID)) DotMatrixDisplay_320 (.clk(clk), .rst(rst), .en_y(wire_6[0:0]), .en_x(wire_33[0:0]), .color_info(wire_6), .pixel_info(wire_33));
  TC_DotMatrixDisplay # (.UUID(64'd832151852570184286 ^ UUID)) DotMatrixDisplay_321 (.clk(clk), .rst(rst), .en_y(wire_67[0:0]), .en_x(wire_33[0:0]), .color_info(wire_67), .pixel_info(wire_33));
  TC_DotMatrixDisplay # (.UUID(64'd2309107926391717062 ^ UUID)) DotMatrixDisplay_322 (.clk(clk), .rst(rst), .en_y(wire_44[0:0]), .en_x(wire_33[0:0]), .color_info(wire_44), .pixel_info(wire_33));
  TC_DotMatrixDisplay # (.UUID(64'd2029970277883025859 ^ UUID)) DotMatrixDisplay_323 (.clk(clk), .rst(rst), .en_y(wire_49[0:0]), .en_x(wire_33[0:0]), .color_info(wire_49), .pixel_info(wire_33));
  TC_DotMatrixDisplay # (.UUID(64'd3674542798305153258 ^ UUID)) DotMatrixDisplay_324 (.clk(clk), .rst(rst), .en_y(wire_71[0:0]), .en_x(wire_33[0:0]), .color_info(wire_71), .pixel_info(wire_33));
  TC_DotMatrixDisplay # (.UUID(64'd1729966332007768227 ^ UUID)) DotMatrixDisplay_325 (.clk(clk), .rst(rst), .en_y(wire_1[0:0]), .en_x(wire_33[0:0]), .color_info(wire_1), .pixel_info(wire_33));
  TC_DotMatrixDisplay # (.UUID(64'd2058241069799366782 ^ UUID)) DotMatrixDisplay_326 (.clk(clk), .rst(rst), .en_y(wire_111[0:0]), .en_x(wire_2[0:0]), .color_info(wire_111), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd2865219518751976828 ^ UUID)) DotMatrixDisplay_327 (.clk(clk), .rst(rst), .en_y(wire_6[0:0]), .en_x(wire_2[0:0]), .color_info(wire_6), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd681129630336150553 ^ UUID)) DotMatrixDisplay_328 (.clk(clk), .rst(rst), .en_y(wire_67[0:0]), .en_x(wire_2[0:0]), .color_info(wire_67), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd1663386889814949500 ^ UUID)) DotMatrixDisplay_329 (.clk(clk), .rst(rst), .en_y(wire_44[0:0]), .en_x(wire_2[0:0]), .color_info(wire_44), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd808553748226111476 ^ UUID)) DotMatrixDisplay_330 (.clk(clk), .rst(rst), .en_y(wire_49[0:0]), .en_x(wire_2[0:0]), .color_info(wire_49), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd746415903002257927 ^ UUID)) DotMatrixDisplay_331 (.clk(clk), .rst(rst), .en_y(wire_71[0:0]), .en_x(wire_2[0:0]), .color_info(wire_71), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd3099060427635950973 ^ UUID)) DotMatrixDisplay_332 (.clk(clk), .rst(rst), .en_y(wire_1[0:0]), .en_x(wire_2[0:0]), .color_info(wire_1), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd846411162372763518 ^ UUID)) DotMatrixDisplay_333 (.clk(clk), .rst(rst), .en_y(wire_111[0:0]), .en_x(wire_47[0:0]), .color_info(wire_111), .pixel_info(wire_47));
  TC_DotMatrixDisplay # (.UUID(64'd2532781995045748377 ^ UUID)) DotMatrixDisplay_334 (.clk(clk), .rst(rst), .en_y(wire_6[0:0]), .en_x(wire_47[0:0]), .color_info(wire_6), .pixel_info(wire_47));
  TC_DotMatrixDisplay # (.UUID(64'd3113666185269458156 ^ UUID)) DotMatrixDisplay_335 (.clk(clk), .rst(rst), .en_y(wire_67[0:0]), .en_x(wire_47[0:0]), .color_info(wire_67), .pixel_info(wire_47));
  TC_DotMatrixDisplay # (.UUID(64'd1236596962882655087 ^ UUID)) DotMatrixDisplay_336 (.clk(clk), .rst(rst), .en_y(wire_44[0:0]), .en_x(wire_47[0:0]), .color_info(wire_44), .pixel_info(wire_47));
  TC_DotMatrixDisplay # (.UUID(64'd4057859383988115461 ^ UUID)) DotMatrixDisplay_337 (.clk(clk), .rst(rst), .en_y(wire_49[0:0]), .en_x(wire_47[0:0]), .color_info(wire_49), .pixel_info(wire_47));
  TC_DotMatrixDisplay # (.UUID(64'd4152225100340615024 ^ UUID)) DotMatrixDisplay_338 (.clk(clk), .rst(rst), .en_y(wire_71[0:0]), .en_x(wire_47[0:0]), .color_info(wire_71), .pixel_info(wire_47));
  TC_DotMatrixDisplay # (.UUID(64'd75066901314019913 ^ UUID)) DotMatrixDisplay_339 (.clk(clk), .rst(rst), .en_y(wire_1[0:0]), .en_x(wire_47[0:0]), .color_info(wire_1), .pixel_info(wire_47));
  TC_DotMatrixDisplay # (.UUID(64'd1809333238917923262 ^ UUID)) DotMatrixDisplay_340 (.clk(clk), .rst(rst), .en_y(wire_6[0:0]), .en_x(wire_31[0:0]), .color_info(wire_6), .pixel_info(wire_31));
  TC_DotMatrixDisplay # (.UUID(64'd39799894064791209 ^ UUID)) DotMatrixDisplay_341 (.clk(clk), .rst(rst), .en_y(wire_67[0:0]), .en_x(wire_31[0:0]), .color_info(wire_67), .pixel_info(wire_31));
  TC_DotMatrixDisplay # (.UUID(64'd443119398778932317 ^ UUID)) DotMatrixDisplay_342 (.clk(clk), .rst(rst), .en_y(wire_44[0:0]), .en_x(wire_31[0:0]), .color_info(wire_44), .pixel_info(wire_31));
  TC_DotMatrixDisplay # (.UUID(64'd3478055426087783047 ^ UUID)) DotMatrixDisplay_343 (.clk(clk), .rst(rst), .en_y(wire_49[0:0]), .en_x(wire_31[0:0]), .color_info(wire_49), .pixel_info(wire_31));
  TC_DotMatrixDisplay # (.UUID(64'd4249516278004530400 ^ UUID)) DotMatrixDisplay_344 (.clk(clk), .rst(rst), .en_y(wire_71[0:0]), .en_x(wire_31[0:0]), .color_info(wire_71), .pixel_info(wire_31));
  TC_DotMatrixDisplay # (.UUID(64'd852854628801789988 ^ UUID)) DotMatrixDisplay_345 (.clk(clk), .rst(rst), .en_y(wire_1[0:0]), .en_x(wire_31[0:0]), .color_info(wire_1), .pixel_info(wire_31));
  TC_DotMatrixDisplay # (.UUID(64'd862426812403186251 ^ UUID)) DotMatrixDisplay_346 (.clk(clk), .rst(rst), .en_y(wire_102[0:0]), .en_x(wire_38[0:0]), .color_info(wire_102), .pixel_info(wire_38));
  TC_DotMatrixDisplay # (.UUID(64'd1175583068235871674 ^ UUID)) DotMatrixDisplay_347 (.clk(clk), .rst(rst), .en_y(wire_113[0:0]), .en_x(wire_38[0:0]), .color_info(wire_113), .pixel_info(wire_38));
  TC_DotMatrixDisplay # (.UUID(64'd1968956125087856272 ^ UUID)) DotMatrixDisplay_348 (.clk(clk), .rst(rst), .en_y(wire_42[0:0]), .en_x(wire_38[0:0]), .color_info(wire_42), .pixel_info(wire_38));
  TC_DotMatrixDisplay # (.UUID(64'd3695429995316965409 ^ UUID)) DotMatrixDisplay_349 (.clk(clk), .rst(rst), .en_y(wire_13[0:0]), .en_x(wire_38[0:0]), .color_info(wire_13), .pixel_info(wire_38));
  TC_DotMatrixDisplay # (.UUID(64'd4426057052600395840 ^ UUID)) DotMatrixDisplay_350 (.clk(clk), .rst(rst), .en_y(wire_92[0:0]), .en_x(wire_38[0:0]), .color_info(wire_92), .pixel_info(wire_38));
  TC_DotMatrixDisplay # (.UUID(64'd1853709868605748700 ^ UUID)) DotMatrixDisplay_351 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_38[0:0]), .color_info(wire_22), .pixel_info(wire_38));
  TC_DotMatrixDisplay # (.UUID(64'd187853449542936450 ^ UUID)) DotMatrixDisplay_352 (.clk(clk), .rst(rst), .en_y(wire_45[0:0]), .en_x(wire_38[0:0]), .color_info(wire_45), .pixel_info(wire_38));
  TC_DotMatrixDisplay # (.UUID(64'd3631399041058968075 ^ UUID)) DotMatrixDisplay_353 (.clk(clk), .rst(rst), .en_y(wire_102[0:0]), .en_x(wire_46[0:0]), .color_info(wire_102), .pixel_info(wire_46));
  TC_DotMatrixDisplay # (.UUID(64'd2290748114189702634 ^ UUID)) DotMatrixDisplay_354 (.clk(clk), .rst(rst), .en_y(wire_113[0:0]), .en_x(wire_46[0:0]), .color_info(wire_113), .pixel_info(wire_46));
  TC_DotMatrixDisplay # (.UUID(64'd1110462014575427719 ^ UUID)) DotMatrixDisplay_355 (.clk(clk), .rst(rst), .en_y(wire_42[0:0]), .en_x(wire_46[0:0]), .color_info(wire_42), .pixel_info(wire_46));
  TC_DotMatrixDisplay # (.UUID(64'd729262243527148738 ^ UUID)) DotMatrixDisplay_356 (.clk(clk), .rst(rst), .en_y(wire_13[0:0]), .en_x(wire_46[0:0]), .color_info(wire_13), .pixel_info(wire_46));
  TC_DotMatrixDisplay # (.UUID(64'd420011481994543514 ^ UUID)) DotMatrixDisplay_357 (.clk(clk), .rst(rst), .en_y(wire_92[0:0]), .en_x(wire_46[0:0]), .color_info(wire_92), .pixel_info(wire_46));
  TC_DotMatrixDisplay # (.UUID(64'd208686899025254723 ^ UUID)) DotMatrixDisplay_358 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_46[0:0]), .color_info(wire_22), .pixel_info(wire_46));
  TC_DotMatrixDisplay # (.UUID(64'd945440528868386831 ^ UUID)) DotMatrixDisplay_359 (.clk(clk), .rst(rst), .en_y(wire_45[0:0]), .en_x(wire_46[0:0]), .color_info(wire_45), .pixel_info(wire_46));
  TC_DotMatrixDisplay # (.UUID(64'd3672409790152176134 ^ UUID)) DotMatrixDisplay_360 (.clk(clk), .rst(rst), .en_y(wire_102[0:0]), .en_x(wire_16[0:0]), .color_info(wire_102), .pixel_info(wire_16));
  TC_DotMatrixDisplay # (.UUID(64'd50498104854955748 ^ UUID)) DotMatrixDisplay_361 (.clk(clk), .rst(rst), .en_y(wire_113[0:0]), .en_x(wire_16[0:0]), .color_info(wire_113), .pixel_info(wire_16));
  TC_DotMatrixDisplay # (.UUID(64'd3066938425878385737 ^ UUID)) DotMatrixDisplay_362 (.clk(clk), .rst(rst), .en_y(wire_42[0:0]), .en_x(wire_16[0:0]), .color_info(wire_42), .pixel_info(wire_16));
  TC_DotMatrixDisplay # (.UUID(64'd452900325122628714 ^ UUID)) DotMatrixDisplay_363 (.clk(clk), .rst(rst), .en_y(wire_13[0:0]), .en_x(wire_16[0:0]), .color_info(wire_13), .pixel_info(wire_16));
  TC_DotMatrixDisplay # (.UUID(64'd1312371312578132690 ^ UUID)) DotMatrixDisplay_364 (.clk(clk), .rst(rst), .en_y(wire_92[0:0]), .en_x(wire_16[0:0]), .color_info(wire_92), .pixel_info(wire_16));
  TC_DotMatrixDisplay # (.UUID(64'd409370946847448641 ^ UUID)) DotMatrixDisplay_365 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_16[0:0]), .color_info(wire_22), .pixel_info(wire_16));
  TC_DotMatrixDisplay # (.UUID(64'd1714045909843845775 ^ UUID)) DotMatrixDisplay_366 (.clk(clk), .rst(rst), .en_y(wire_45[0:0]), .en_x(wire_16[0:0]), .color_info(wire_45), .pixel_info(wire_16));
  TC_DotMatrixDisplay # (.UUID(64'd582973553920656968 ^ UUID)) DotMatrixDisplay_367 (.clk(clk), .rst(rst), .en_y(wire_102[0:0]), .en_x(wire_11[0:0]), .color_info(wire_102), .pixel_info(wire_11));
  TC_DotMatrixDisplay # (.UUID(64'd1091068617740911605 ^ UUID)) DotMatrixDisplay_368 (.clk(clk), .rst(rst), .en_y(wire_113[0:0]), .en_x(wire_11[0:0]), .color_info(wire_113), .pixel_info(wire_11));
  TC_DotMatrixDisplay # (.UUID(64'd2090984655901458436 ^ UUID)) DotMatrixDisplay_369 (.clk(clk), .rst(rst), .en_y(wire_42[0:0]), .en_x(wire_11[0:0]), .color_info(wire_42), .pixel_info(wire_11));
  TC_DotMatrixDisplay # (.UUID(64'd1567590639541441330 ^ UUID)) DotMatrixDisplay_370 (.clk(clk), .rst(rst), .en_y(wire_13[0:0]), .en_x(wire_11[0:0]), .color_info(wire_13), .pixel_info(wire_11));
  TC_DotMatrixDisplay # (.UUID(64'd4551077945493198585 ^ UUID)) DotMatrixDisplay_371 (.clk(clk), .rst(rst), .en_y(wire_92[0:0]), .en_x(wire_11[0:0]), .color_info(wire_92), .pixel_info(wire_11));
  TC_DotMatrixDisplay # (.UUID(64'd4550724431840064912 ^ UUID)) DotMatrixDisplay_372 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_11[0:0]), .color_info(wire_22), .pixel_info(wire_11));
  TC_DotMatrixDisplay # (.UUID(64'd965320783751459911 ^ UUID)) DotMatrixDisplay_373 (.clk(clk), .rst(rst), .en_y(wire_45[0:0]), .en_x(wire_11[0:0]), .color_info(wire_45), .pixel_info(wire_11));
  TC_DotMatrixDisplay # (.UUID(64'd4051602518287011043 ^ UUID)) DotMatrixDisplay_374 (.clk(clk), .rst(rst), .en_y(wire_102[0:0]), .en_x(wire_65[0:0]), .color_info(wire_102), .pixel_info(wire_65));
  TC_DotMatrixDisplay # (.UUID(64'd2296309809473862596 ^ UUID)) DotMatrixDisplay_375 (.clk(clk), .rst(rst), .en_y(wire_113[0:0]), .en_x(wire_65[0:0]), .color_info(wire_113), .pixel_info(wire_65));
  TC_DotMatrixDisplay # (.UUID(64'd1788635125803614051 ^ UUID)) DotMatrixDisplay_376 (.clk(clk), .rst(rst), .en_y(wire_42[0:0]), .en_x(wire_65[0:0]), .color_info(wire_42), .pixel_info(wire_65));
  TC_DotMatrixDisplay # (.UUID(64'd122586930798985372 ^ UUID)) DotMatrixDisplay_377 (.clk(clk), .rst(rst), .en_y(wire_13[0:0]), .en_x(wire_65[0:0]), .color_info(wire_13), .pixel_info(wire_65));
  TC_DotMatrixDisplay # (.UUID(64'd3150935394061164609 ^ UUID)) DotMatrixDisplay_378 (.clk(clk), .rst(rst), .en_y(wire_92[0:0]), .en_x(wire_65[0:0]), .color_info(wire_92), .pixel_info(wire_65));
  TC_DotMatrixDisplay # (.UUID(64'd695681827614291978 ^ UUID)) DotMatrixDisplay_379 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_65[0:0]), .color_info(wire_22), .pixel_info(wire_65));
  TC_DotMatrixDisplay # (.UUID(64'd4222155341837459308 ^ UUID)) DotMatrixDisplay_380 (.clk(clk), .rst(rst), .en_y(wire_45[0:0]), .en_x(wire_65[0:0]), .color_info(wire_45), .pixel_info(wire_65));
  TC_DotMatrixDisplay # (.UUID(64'd4287440396605129792 ^ UUID)) DotMatrixDisplay_381 (.clk(clk), .rst(rst), .en_y(wire_102[0:0]), .en_x(wire_7[0:0]), .color_info(wire_102), .pixel_info(wire_7));
  TC_DotMatrixDisplay # (.UUID(64'd2535731812463731870 ^ UUID)) DotMatrixDisplay_382 (.clk(clk), .rst(rst), .en_y(wire_113[0:0]), .en_x(wire_7[0:0]), .color_info(wire_113), .pixel_info(wire_7));
  TC_DotMatrixDisplay # (.UUID(64'd3795774870147768231 ^ UUID)) DotMatrixDisplay_383 (.clk(clk), .rst(rst), .en_y(wire_42[0:0]), .en_x(wire_7[0:0]), .color_info(wire_42), .pixel_info(wire_7));
  TC_DotMatrixDisplay # (.UUID(64'd4186020613379327615 ^ UUID)) DotMatrixDisplay_384 (.clk(clk), .rst(rst), .en_y(wire_13[0:0]), .en_x(wire_7[0:0]), .color_info(wire_13), .pixel_info(wire_7));
  TC_DotMatrixDisplay # (.UUID(64'd3654035419741017261 ^ UUID)) DotMatrixDisplay_385 (.clk(clk), .rst(rst), .en_y(wire_92[0:0]), .en_x(wire_7[0:0]), .color_info(wire_92), .pixel_info(wire_7));
  TC_DotMatrixDisplay # (.UUID(64'd3593055696864145732 ^ UUID)) DotMatrixDisplay_386 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_7[0:0]), .color_info(wire_22), .pixel_info(wire_7));
  TC_DotMatrixDisplay # (.UUID(64'd4051058533280774412 ^ UUID)) DotMatrixDisplay_387 (.clk(clk), .rst(rst), .en_y(wire_45[0:0]), .en_x(wire_7[0:0]), .color_info(wire_45), .pixel_info(wire_7));
  TC_DotMatrixDisplay # (.UUID(64'd230567006613948312 ^ UUID)) DotMatrixDisplay_388 (.clk(clk), .rst(rst), .en_y(wire_92[0:0]), .en_x(wire_52[0:0]), .color_info(wire_92), .pixel_info(wire_52));
  TC_DotMatrixDisplay # (.UUID(64'd3674494280367613976 ^ UUID)) DotMatrixDisplay_389 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_52[0:0]), .color_info(wire_22), .pixel_info(wire_52));
  TC_DotMatrixDisplay # (.UUID(64'd1902890806744483172 ^ UUID)) DotMatrixDisplay_390 (.clk(clk), .rst(rst), .en_y(wire_45[0:0]), .en_x(wire_52[0:0]), .color_info(wire_45), .pixel_info(wire_52));
  TC_DotMatrixDisplay # (.UUID(64'd3058636886864204816 ^ UUID)) DotMatrixDisplay_391 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_41[0:0]), .color_info(wire_22), .pixel_info(wire_41));
  TC_DotMatrixDisplay # (.UUID(64'd3302876998549722765 ^ UUID)) DotMatrixDisplay_392 (.clk(clk), .rst(rst), .en_y(wire_45[0:0]), .en_x(wire_41[0:0]), .color_info(wire_45), .pixel_info(wire_41));
  TC_DotMatrixDisplay # (.UUID(64'd164050661385911247 ^ UUID)) DotMatrixDisplay_393 (.clk(clk), .rst(rst), .en_y(wire_102[0:0]), .en_x(wire_59[0:0]), .color_info(wire_102), .pixel_info(wire_59));
  TC_DotMatrixDisplay # (.UUID(64'd2211666196312108003 ^ UUID)) DotMatrixDisplay_394 (.clk(clk), .rst(rst), .en_y(wire_113[0:0]), .en_x(wire_59[0:0]), .color_info(wire_113), .pixel_info(wire_59));
  TC_DotMatrixDisplay # (.UUID(64'd1720566550546644761 ^ UUID)) DotMatrixDisplay_395 (.clk(clk), .rst(rst), .en_y(wire_42[0:0]), .en_x(wire_59[0:0]), .color_info(wire_42), .pixel_info(wire_59));
  TC_DotMatrixDisplay # (.UUID(64'd963115573635329400 ^ UUID)) DotMatrixDisplay_396 (.clk(clk), .rst(rst), .en_y(wire_13[0:0]), .en_x(wire_59[0:0]), .color_info(wire_13), .pixel_info(wire_59));
  TC_DotMatrixDisplay # (.UUID(64'd1587438248241797071 ^ UUID)) DotMatrixDisplay_397 (.clk(clk), .rst(rst), .en_y(wire_92[0:0]), .en_x(wire_59[0:0]), .color_info(wire_92), .pixel_info(wire_59));
  TC_DotMatrixDisplay # (.UUID(64'd2284191432046994452 ^ UUID)) DotMatrixDisplay_398 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_59[0:0]), .color_info(wire_22), .pixel_info(wire_59));
  TC_DotMatrixDisplay # (.UUID(64'd2321204376582881813 ^ UUID)) DotMatrixDisplay_399 (.clk(clk), .rst(rst), .en_y(wire_45[0:0]), .en_x(wire_59[0:0]), .color_info(wire_45), .pixel_info(wire_59));
  TC_DotMatrixDisplay # (.UUID(64'd3791930441930289359 ^ UUID)) DotMatrixDisplay_400 (.clk(clk), .rst(rst), .en_y(wire_102[0:0]), .en_x(wire_30[0:0]), .color_info(wire_102), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd2521732661635123702 ^ UUID)) DotMatrixDisplay_401 (.clk(clk), .rst(rst), .en_y(wire_113[0:0]), .en_x(wire_30[0:0]), .color_info(wire_113), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd4052107426107744403 ^ UUID)) DotMatrixDisplay_402 (.clk(clk), .rst(rst), .en_y(wire_42[0:0]), .en_x(wire_30[0:0]), .color_info(wire_42), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd3969114452687428160 ^ UUID)) DotMatrixDisplay_403 (.clk(clk), .rst(rst), .en_y(wire_13[0:0]), .en_x(wire_30[0:0]), .color_info(wire_13), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd2757689911680787592 ^ UUID)) DotMatrixDisplay_404 (.clk(clk), .rst(rst), .en_y(wire_92[0:0]), .en_x(wire_30[0:0]), .color_info(wire_92), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd1728098641799782145 ^ UUID)) DotMatrixDisplay_405 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_30[0:0]), .color_info(wire_22), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd663883931804341073 ^ UUID)) DotMatrixDisplay_406 (.clk(clk), .rst(rst), .en_y(wire_45[0:0]), .en_x(wire_30[0:0]), .color_info(wire_45), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd1125836511926786919 ^ UUID)) DotMatrixDisplay_407 (.clk(clk), .rst(rst), .en_y(wire_102[0:0]), .en_x(wire_57[0:0]), .color_info(wire_102), .pixel_info(wire_57));
  TC_DotMatrixDisplay # (.UUID(64'd1635922883591559242 ^ UUID)) DotMatrixDisplay_408 (.clk(clk), .rst(rst), .en_y(wire_113[0:0]), .en_x(wire_57[0:0]), .color_info(wire_113), .pixel_info(wire_57));
  TC_DotMatrixDisplay # (.UUID(64'd1549700521013509780 ^ UUID)) DotMatrixDisplay_409 (.clk(clk), .rst(rst), .en_y(wire_42[0:0]), .en_x(wire_57[0:0]), .color_info(wire_42), .pixel_info(wire_57));
  TC_DotMatrixDisplay # (.UUID(64'd1126192879190487974 ^ UUID)) DotMatrixDisplay_410 (.clk(clk), .rst(rst), .en_y(wire_13[0:0]), .en_x(wire_57[0:0]), .color_info(wire_13), .pixel_info(wire_57));
  TC_DotMatrixDisplay # (.UUID(64'd539245102989418868 ^ UUID)) DotMatrixDisplay_411 (.clk(clk), .rst(rst), .en_y(wire_92[0:0]), .en_x(wire_57[0:0]), .color_info(wire_92), .pixel_info(wire_57));
  TC_DotMatrixDisplay # (.UUID(64'd1581959596343711711 ^ UUID)) DotMatrixDisplay_412 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_57[0:0]), .color_info(wire_22), .pixel_info(wire_57));
  TC_DotMatrixDisplay # (.UUID(64'd64401492364826964 ^ UUID)) DotMatrixDisplay_413 (.clk(clk), .rst(rst), .en_y(wire_45[0:0]), .en_x(wire_57[0:0]), .color_info(wire_45), .pixel_info(wire_57));
  TC_DotMatrixDisplay # (.UUID(64'd4525768993628488402 ^ UUID)) DotMatrixDisplay_414 (.clk(clk), .rst(rst), .en_y(wire_102[0:0]), .en_x(wire_33[0:0]), .color_info(wire_102), .pixel_info(wire_33));
  TC_DotMatrixDisplay # (.UUID(64'd2115176533976111260 ^ UUID)) DotMatrixDisplay_415 (.clk(clk), .rst(rst), .en_y(wire_113[0:0]), .en_x(wire_33[0:0]), .color_info(wire_113), .pixel_info(wire_33));
  TC_DotMatrixDisplay # (.UUID(64'd909317690909131686 ^ UUID)) DotMatrixDisplay_416 (.clk(clk), .rst(rst), .en_y(wire_42[0:0]), .en_x(wire_33[0:0]), .color_info(wire_42), .pixel_info(wire_33));
  TC_DotMatrixDisplay # (.UUID(64'd3073197554694154441 ^ UUID)) DotMatrixDisplay_417 (.clk(clk), .rst(rst), .en_y(wire_13[0:0]), .en_x(wire_33[0:0]), .color_info(wire_13), .pixel_info(wire_33));
  TC_DotMatrixDisplay # (.UUID(64'd845952556993319905 ^ UUID)) DotMatrixDisplay_418 (.clk(clk), .rst(rst), .en_y(wire_92[0:0]), .en_x(wire_33[0:0]), .color_info(wire_92), .pixel_info(wire_33));
  TC_DotMatrixDisplay # (.UUID(64'd2342725993517367987 ^ UUID)) DotMatrixDisplay_419 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_33[0:0]), .color_info(wire_22), .pixel_info(wire_33));
  TC_DotMatrixDisplay # (.UUID(64'd2090786563299024876 ^ UUID)) DotMatrixDisplay_420 (.clk(clk), .rst(rst), .en_y(wire_45[0:0]), .en_x(wire_33[0:0]), .color_info(wire_45), .pixel_info(wire_33));
  TC_DotMatrixDisplay # (.UUID(64'd308814793204862390 ^ UUID)) DotMatrixDisplay_421 (.clk(clk), .rst(rst), .en_y(wire_102[0:0]), .en_x(wire_2[0:0]), .color_info(wire_102), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd756518983919304125 ^ UUID)) DotMatrixDisplay_422 (.clk(clk), .rst(rst), .en_y(wire_113[0:0]), .en_x(wire_2[0:0]), .color_info(wire_113), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd868029179401946150 ^ UUID)) DotMatrixDisplay_423 (.clk(clk), .rst(rst), .en_y(wire_42[0:0]), .en_x(wire_2[0:0]), .color_info(wire_42), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd3086534555144355480 ^ UUID)) DotMatrixDisplay_424 (.clk(clk), .rst(rst), .en_y(wire_13[0:0]), .en_x(wire_2[0:0]), .color_info(wire_13), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd2543873466149892510 ^ UUID)) DotMatrixDisplay_425 (.clk(clk), .rst(rst), .en_y(wire_92[0:0]), .en_x(wire_2[0:0]), .color_info(wire_92), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd1263466635050190748 ^ UUID)) DotMatrixDisplay_426 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_2[0:0]), .color_info(wire_22), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd1058264461621773172 ^ UUID)) DotMatrixDisplay_427 (.clk(clk), .rst(rst), .en_y(wire_45[0:0]), .en_x(wire_2[0:0]), .color_info(wire_45), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd3633660340223074985 ^ UUID)) DotMatrixDisplay_428 (.clk(clk), .rst(rst), .en_y(wire_102[0:0]), .en_x(wire_47[0:0]), .color_info(wire_102), .pixel_info(wire_47));
  TC_DotMatrixDisplay # (.UUID(64'd3433076540254304157 ^ UUID)) DotMatrixDisplay_429 (.clk(clk), .rst(rst), .en_y(wire_113[0:0]), .en_x(wire_47[0:0]), .color_info(wire_113), .pixel_info(wire_47));
  TC_DotMatrixDisplay # (.UUID(64'd4203607823351378081 ^ UUID)) DotMatrixDisplay_430 (.clk(clk), .rst(rst), .en_y(wire_42[0:0]), .en_x(wire_47[0:0]), .color_info(wire_42), .pixel_info(wire_47));
  TC_DotMatrixDisplay # (.UUID(64'd3632131432567039130 ^ UUID)) DotMatrixDisplay_431 (.clk(clk), .rst(rst), .en_y(wire_13[0:0]), .en_x(wire_47[0:0]), .color_info(wire_13), .pixel_info(wire_47));
  TC_DotMatrixDisplay # (.UUID(64'd453714807272017425 ^ UUID)) DotMatrixDisplay_432 (.clk(clk), .rst(rst), .en_y(wire_92[0:0]), .en_x(wire_47[0:0]), .color_info(wire_92), .pixel_info(wire_47));
  TC_DotMatrixDisplay # (.UUID(64'd3278495577680984269 ^ UUID)) DotMatrixDisplay_433 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_47[0:0]), .color_info(wire_22), .pixel_info(wire_47));
  TC_DotMatrixDisplay # (.UUID(64'd1319574741952347969 ^ UUID)) DotMatrixDisplay_434 (.clk(clk), .rst(rst), .en_y(wire_45[0:0]), .en_x(wire_47[0:0]), .color_info(wire_45), .pixel_info(wire_47));
  TC_DotMatrixDisplay # (.UUID(64'd1802800560535904000 ^ UUID)) DotMatrixDisplay_435 (.clk(clk), .rst(rst), .en_y(wire_102[0:0]), .en_x(wire_31[0:0]), .color_info(wire_102), .pixel_info(wire_31));
  TC_DotMatrixDisplay # (.UUID(64'd3155257920911904589 ^ UUID)) DotMatrixDisplay_436 (.clk(clk), .rst(rst), .en_y(wire_113[0:0]), .en_x(wire_31[0:0]), .color_info(wire_113), .pixel_info(wire_31));
  TC_DotMatrixDisplay # (.UUID(64'd2312916404027271402 ^ UUID)) DotMatrixDisplay_437 (.clk(clk), .rst(rst), .en_y(wire_42[0:0]), .en_x(wire_31[0:0]), .color_info(wire_42), .pixel_info(wire_31));
  TC_DotMatrixDisplay # (.UUID(64'd770501697257851765 ^ UUID)) DotMatrixDisplay_438 (.clk(clk), .rst(rst), .en_y(wire_13[0:0]), .en_x(wire_31[0:0]), .color_info(wire_13), .pixel_info(wire_31));
  TC_DotMatrixDisplay # (.UUID(64'd3136109271020180467 ^ UUID)) DotMatrixDisplay_439 (.clk(clk), .rst(rst), .en_y(wire_92[0:0]), .en_x(wire_31[0:0]), .color_info(wire_92), .pixel_info(wire_31));
  TC_DotMatrixDisplay # (.UUID(64'd738865139799679064 ^ UUID)) DotMatrixDisplay_440 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_31[0:0]), .color_info(wire_22), .pixel_info(wire_31));
  TC_DotMatrixDisplay # (.UUID(64'd239226686861837210 ^ UUID)) DotMatrixDisplay_441 (.clk(clk), .rst(rst), .en_y(wire_45[0:0]), .en_x(wire_31[0:0]), .color_info(wire_45), .pixel_info(wire_31));
  TC_DotMatrixDisplay # (.UUID(64'd1710146568569270280 ^ UUID)) DotMatrixDisplay_442 (.clk(clk), .rst(rst), .en_y(wire_53[0:0]), .en_x(wire_38[0:0]), .color_info(wire_53), .pixel_info(wire_38));
  TC_DotMatrixDisplay # (.UUID(64'd1892066800965434951 ^ UUID)) DotMatrixDisplay_443 (.clk(clk), .rst(rst), .en_y(wire_66[0:0]), .en_x(wire_38[0:0]), .color_info(wire_66), .pixel_info(wire_38));
  TC_DotMatrixDisplay # (.UUID(64'd2768061308888516295 ^ UUID)) DotMatrixDisplay_444 (.clk(clk), .rst(rst), .en_y(wire_105[0:0]), .en_x(wire_38[0:0]), .color_info(wire_105), .pixel_info(wire_38));
  TC_DotMatrixDisplay # (.UUID(64'd3011302873972680241 ^ UUID)) DotMatrixDisplay_445 (.clk(clk), .rst(rst), .en_y(wire_40[0:0]), .en_x(wire_38[0:0]), .color_info(wire_40), .pixel_info(wire_38));
  TC_DotMatrixDisplay # (.UUID(64'd4064114457568423260 ^ UUID)) DotMatrixDisplay_446 (.clk(clk), .rst(rst), .en_y(wire_69[0:0]), .en_x(wire_38[0:0]), .color_info(wire_69), .pixel_info(wire_38));
  TC_DotMatrixDisplay # (.UUID(64'd2949345132651038803 ^ UUID)) DotMatrixDisplay_447 (.clk(clk), .rst(rst), .en_y(wire_17[0:0]), .en_x(wire_38[0:0]), .color_info(wire_17), .pixel_info(wire_38));
  TC_DotMatrixDisplay # (.UUID(64'd1757104896198618793 ^ UUID)) DotMatrixDisplay_448 (.clk(clk), .rst(rst), .en_y(wire_20[0:0]), .en_x(wire_38[0:0]), .color_info(wire_20), .pixel_info(wire_38));
  TC_DotMatrixDisplay # (.UUID(64'd699790011527599470 ^ UUID)) DotMatrixDisplay_449 (.clk(clk), .rst(rst), .en_y(wire_53[0:0]), .en_x(wire_46[0:0]), .color_info(wire_53), .pixel_info(wire_46));
  TC_DotMatrixDisplay # (.UUID(64'd4559640237467913593 ^ UUID)) DotMatrixDisplay_450 (.clk(clk), .rst(rst), .en_y(wire_66[0:0]), .en_x(wire_46[0:0]), .color_info(wire_66), .pixel_info(wire_46));
  TC_DotMatrixDisplay # (.UUID(64'd3221817849220702119 ^ UUID)) DotMatrixDisplay_451 (.clk(clk), .rst(rst), .en_y(wire_105[0:0]), .en_x(wire_46[0:0]), .color_info(wire_105), .pixel_info(wire_46));
  TC_DotMatrixDisplay # (.UUID(64'd1361453408987900468 ^ UUID)) DotMatrixDisplay_452 (.clk(clk), .rst(rst), .en_y(wire_40[0:0]), .en_x(wire_46[0:0]), .color_info(wire_40), .pixel_info(wire_46));
  TC_DotMatrixDisplay # (.UUID(64'd4119918883605204059 ^ UUID)) DotMatrixDisplay_453 (.clk(clk), .rst(rst), .en_y(wire_69[0:0]), .en_x(wire_46[0:0]), .color_info(wire_69), .pixel_info(wire_46));
  TC_DotMatrixDisplay # (.UUID(64'd2126688544406480223 ^ UUID)) DotMatrixDisplay_454 (.clk(clk), .rst(rst), .en_y(wire_17[0:0]), .en_x(wire_46[0:0]), .color_info(wire_17), .pixel_info(wire_46));
  TC_DotMatrixDisplay # (.UUID(64'd1688371966109459924 ^ UUID)) DotMatrixDisplay_455 (.clk(clk), .rst(rst), .en_y(wire_20[0:0]), .en_x(wire_46[0:0]), .color_info(wire_20), .pixel_info(wire_46));
  TC_DotMatrixDisplay # (.UUID(64'd1405645478306846645 ^ UUID)) DotMatrixDisplay_456 (.clk(clk), .rst(rst), .en_y(wire_53[0:0]), .en_x(wire_16[0:0]), .color_info(wire_53), .pixel_info(wire_16));
  TC_DotMatrixDisplay # (.UUID(64'd3248684792212771849 ^ UUID)) DotMatrixDisplay_457 (.clk(clk), .rst(rst), .en_y(wire_66[0:0]), .en_x(wire_16[0:0]), .color_info(wire_66), .pixel_info(wire_16));
  TC_DotMatrixDisplay # (.UUID(64'd3525457726748371427 ^ UUID)) DotMatrixDisplay_458 (.clk(clk), .rst(rst), .en_y(wire_105[0:0]), .en_x(wire_16[0:0]), .color_info(wire_105), .pixel_info(wire_16));
  TC_DotMatrixDisplay # (.UUID(64'd3211849938453158766 ^ UUID)) DotMatrixDisplay_459 (.clk(clk), .rst(rst), .en_y(wire_40[0:0]), .en_x(wire_16[0:0]), .color_info(wire_40), .pixel_info(wire_16));
  TC_DotMatrixDisplay # (.UUID(64'd4408247672558102839 ^ UUID)) DotMatrixDisplay_460 (.clk(clk), .rst(rst), .en_y(wire_69[0:0]), .en_x(wire_16[0:0]), .color_info(wire_69), .pixel_info(wire_16));
  TC_DotMatrixDisplay # (.UUID(64'd2724859932618838942 ^ UUID)) DotMatrixDisplay_461 (.clk(clk), .rst(rst), .en_y(wire_17[0:0]), .en_x(wire_16[0:0]), .color_info(wire_17), .pixel_info(wire_16));
  TC_DotMatrixDisplay # (.UUID(64'd4423999222896730745 ^ UUID)) DotMatrixDisplay_462 (.clk(clk), .rst(rst), .en_y(wire_20[0:0]), .en_x(wire_16[0:0]), .color_info(wire_20), .pixel_info(wire_16));
  TC_DotMatrixDisplay # (.UUID(64'd410227581406671113 ^ UUID)) DotMatrixDisplay_463 (.clk(clk), .rst(rst), .en_y(wire_53[0:0]), .en_x(wire_11[0:0]), .color_info(wire_53), .pixel_info(wire_11));
  TC_DotMatrixDisplay # (.UUID(64'd1018663185908120475 ^ UUID)) DotMatrixDisplay_464 (.clk(clk), .rst(rst), .en_y(wire_66[0:0]), .en_x(wire_11[0:0]), .color_info(wire_66), .pixel_info(wire_11));
  TC_DotMatrixDisplay # (.UUID(64'd4315192005535331019 ^ UUID)) DotMatrixDisplay_465 (.clk(clk), .rst(rst), .en_y(wire_105[0:0]), .en_x(wire_11[0:0]), .color_info(wire_105), .pixel_info(wire_11));
  TC_DotMatrixDisplay # (.UUID(64'd3858179522860762253 ^ UUID)) DotMatrixDisplay_466 (.clk(clk), .rst(rst), .en_y(wire_40[0:0]), .en_x(wire_11[0:0]), .color_info(wire_40), .pixel_info(wire_11));
  TC_DotMatrixDisplay # (.UUID(64'd2233108556641031856 ^ UUID)) DotMatrixDisplay_467 (.clk(clk), .rst(rst), .en_y(wire_69[0:0]), .en_x(wire_11[0:0]), .color_info(wire_69), .pixel_info(wire_11));
  TC_DotMatrixDisplay # (.UUID(64'd341403828675164188 ^ UUID)) DotMatrixDisplay_468 (.clk(clk), .rst(rst), .en_y(wire_17[0:0]), .en_x(wire_11[0:0]), .color_info(wire_17), .pixel_info(wire_11));
  TC_DotMatrixDisplay # (.UUID(64'd4502986987875139623 ^ UUID)) DotMatrixDisplay_469 (.clk(clk), .rst(rst), .en_y(wire_20[0:0]), .en_x(wire_11[0:0]), .color_info(wire_20), .pixel_info(wire_11));
  TC_DotMatrixDisplay # (.UUID(64'd2472304368392065306 ^ UUID)) DotMatrixDisplay_470 (.clk(clk), .rst(rst), .en_y(wire_53[0:0]), .en_x(wire_65[0:0]), .color_info(wire_53), .pixel_info(wire_65));
  TC_DotMatrixDisplay # (.UUID(64'd388702590735162125 ^ UUID)) DotMatrixDisplay_471 (.clk(clk), .rst(rst), .en_y(wire_66[0:0]), .en_x(wire_65[0:0]), .color_info(wire_66), .pixel_info(wire_65));
  TC_DotMatrixDisplay # (.UUID(64'd4349947969052345094 ^ UUID)) DotMatrixDisplay_472 (.clk(clk), .rst(rst), .en_y(wire_105[0:0]), .en_x(wire_65[0:0]), .color_info(wire_105), .pixel_info(wire_65));
  TC_DotMatrixDisplay # (.UUID(64'd2830186379754490470 ^ UUID)) DotMatrixDisplay_473 (.clk(clk), .rst(rst), .en_y(wire_40[0:0]), .en_x(wire_65[0:0]), .color_info(wire_40), .pixel_info(wire_65));
  TC_DotMatrixDisplay # (.UUID(64'd2751237613574193307 ^ UUID)) DotMatrixDisplay_474 (.clk(clk), .rst(rst), .en_y(wire_69[0:0]), .en_x(wire_65[0:0]), .color_info(wire_69), .pixel_info(wire_65));
  TC_DotMatrixDisplay # (.UUID(64'd2368716884893433047 ^ UUID)) DotMatrixDisplay_475 (.clk(clk), .rst(rst), .en_y(wire_17[0:0]), .en_x(wire_65[0:0]), .color_info(wire_17), .pixel_info(wire_65));
  TC_DotMatrixDisplay # (.UUID(64'd1475085101361714055 ^ UUID)) DotMatrixDisplay_476 (.clk(clk), .rst(rst), .en_y(wire_20[0:0]), .en_x(wire_65[0:0]), .color_info(wire_20), .pixel_info(wire_65));
  TC_DotMatrixDisplay # (.UUID(64'd3103815246634105942 ^ UUID)) DotMatrixDisplay_477 (.clk(clk), .rst(rst), .en_y(wire_53[0:0]), .en_x(wire_7[0:0]), .color_info(wire_53), .pixel_info(wire_7));
  TC_DotMatrixDisplay # (.UUID(64'd1870390980476747323 ^ UUID)) DotMatrixDisplay_478 (.clk(clk), .rst(rst), .en_y(wire_66[0:0]), .en_x(wire_7[0:0]), .color_info(wire_66), .pixel_info(wire_7));
  TC_DotMatrixDisplay # (.UUID(64'd2465358875045855314 ^ UUID)) DotMatrixDisplay_479 (.clk(clk), .rst(rst), .en_y(wire_105[0:0]), .en_x(wire_7[0:0]), .color_info(wire_105), .pixel_info(wire_7));
  TC_DotMatrixDisplay # (.UUID(64'd2617578140411458120 ^ UUID)) DotMatrixDisplay_480 (.clk(clk), .rst(rst), .en_y(wire_40[0:0]), .en_x(wire_7[0:0]), .color_info(wire_40), .pixel_info(wire_7));
  TC_DotMatrixDisplay # (.UUID(64'd2589744481661745670 ^ UUID)) DotMatrixDisplay_481 (.clk(clk), .rst(rst), .en_y(wire_69[0:0]), .en_x(wire_7[0:0]), .color_info(wire_69), .pixel_info(wire_7));
  TC_DotMatrixDisplay # (.UUID(64'd2005384577281396007 ^ UUID)) DotMatrixDisplay_482 (.clk(clk), .rst(rst), .en_y(wire_17[0:0]), .en_x(wire_7[0:0]), .color_info(wire_17), .pixel_info(wire_7));
  TC_DotMatrixDisplay # (.UUID(64'd402546619115129690 ^ UUID)) DotMatrixDisplay_483 (.clk(clk), .rst(rst), .en_y(wire_20[0:0]), .en_x(wire_7[0:0]), .color_info(wire_20), .pixel_info(wire_7));
  TC_DotMatrixDisplay # (.UUID(64'd3742423865784027785 ^ UUID)) DotMatrixDisplay_484 (.clk(clk), .rst(rst), .en_y(wire_53[0:0]), .en_x(wire_52[0:0]), .color_info(wire_53), .pixel_info(wire_52));
  TC_DotMatrixDisplay # (.UUID(64'd5226187604462580 ^ UUID)) DotMatrixDisplay_485 (.clk(clk), .rst(rst), .en_y(wire_66[0:0]), .en_x(wire_52[0:0]), .color_info(wire_66), .pixel_info(wire_52));
  TC_DotMatrixDisplay # (.UUID(64'd3404708907280667073 ^ UUID)) DotMatrixDisplay_486 (.clk(clk), .rst(rst), .en_y(wire_105[0:0]), .en_x(wire_52[0:0]), .color_info(wire_105), .pixel_info(wire_52));
  TC_DotMatrixDisplay # (.UUID(64'd216126835035472207 ^ UUID)) DotMatrixDisplay_487 (.clk(clk), .rst(rst), .en_y(wire_40[0:0]), .en_x(wire_52[0:0]), .color_info(wire_40), .pixel_info(wire_52));
  TC_DotMatrixDisplay # (.UUID(64'd1306148363587124625 ^ UUID)) DotMatrixDisplay_488 (.clk(clk), .rst(rst), .en_y(wire_69[0:0]), .en_x(wire_52[0:0]), .color_info(wire_69), .pixel_info(wire_52));
  TC_DotMatrixDisplay # (.UUID(64'd783780666640220283 ^ UUID)) DotMatrixDisplay_489 (.clk(clk), .rst(rst), .en_y(wire_17[0:0]), .en_x(wire_52[0:0]), .color_info(wire_17), .pixel_info(wire_52));
  TC_DotMatrixDisplay # (.UUID(64'd4532985192935913249 ^ UUID)) DotMatrixDisplay_490 (.clk(clk), .rst(rst), .en_y(wire_20[0:0]), .en_x(wire_52[0:0]), .color_info(wire_20), .pixel_info(wire_52));
  TC_DotMatrixDisplay # (.UUID(64'd1062857310501978557 ^ UUID)) DotMatrixDisplay_491 (.clk(clk), .rst(rst), .en_y(wire_53[0:0]), .en_x(wire_41[0:0]), .color_info(wire_53), .pixel_info(wire_41));
  TC_DotMatrixDisplay # (.UUID(64'd3760687265496207315 ^ UUID)) DotMatrixDisplay_492 (.clk(clk), .rst(rst), .en_y(wire_66[0:0]), .en_x(wire_41[0:0]), .color_info(wire_66), .pixel_info(wire_41));
  TC_DotMatrixDisplay # (.UUID(64'd3937456510983979812 ^ UUID)) DotMatrixDisplay_493 (.clk(clk), .rst(rst), .en_y(wire_105[0:0]), .en_x(wire_41[0:0]), .color_info(wire_105), .pixel_info(wire_41));
  TC_DotMatrixDisplay # (.UUID(64'd3373365589932917652 ^ UUID)) DotMatrixDisplay_494 (.clk(clk), .rst(rst), .en_y(wire_40[0:0]), .en_x(wire_41[0:0]), .color_info(wire_40), .pixel_info(wire_41));
  TC_DotMatrixDisplay # (.UUID(64'd1988819457438404312 ^ UUID)) DotMatrixDisplay_495 (.clk(clk), .rst(rst), .en_y(wire_69[0:0]), .en_x(wire_41[0:0]), .color_info(wire_69), .pixel_info(wire_41));
  TC_DotMatrixDisplay # (.UUID(64'd3660006191238004380 ^ UUID)) DotMatrixDisplay_496 (.clk(clk), .rst(rst), .en_y(wire_17[0:0]), .en_x(wire_41[0:0]), .color_info(wire_17), .pixel_info(wire_41));
  TC_DotMatrixDisplay # (.UUID(64'd4120680415267466967 ^ UUID)) DotMatrixDisplay_497 (.clk(clk), .rst(rst), .en_y(wire_20[0:0]), .en_x(wire_41[0:0]), .color_info(wire_20), .pixel_info(wire_41));
  TC_DotMatrixDisplay # (.UUID(64'd1966982712986781527 ^ UUID)) DotMatrixDisplay_498 (.clk(clk), .rst(rst), .en_y(wire_53[0:0]), .en_x(wire_59[0:0]), .color_info(wire_53), .pixel_info(wire_59));
  TC_DotMatrixDisplay # (.UUID(64'd2816617433896888837 ^ UUID)) DotMatrixDisplay_499 (.clk(clk), .rst(rst), .en_y(wire_66[0:0]), .en_x(wire_59[0:0]), .color_info(wire_66), .pixel_info(wire_59));
  TC_DotMatrixDisplay # (.UUID(64'd2473485147585956800 ^ UUID)) DotMatrixDisplay_500 (.clk(clk), .rst(rst), .en_y(wire_105[0:0]), .en_x(wire_59[0:0]), .color_info(wire_105), .pixel_info(wire_59));
  TC_DotMatrixDisplay # (.UUID(64'd269647066566553933 ^ UUID)) DotMatrixDisplay_501 (.clk(clk), .rst(rst), .en_y(wire_40[0:0]), .en_x(wire_59[0:0]), .color_info(wire_40), .pixel_info(wire_59));
  TC_DotMatrixDisplay # (.UUID(64'd919624889098312256 ^ UUID)) DotMatrixDisplay_502 (.clk(clk), .rst(rst), .en_y(wire_69[0:0]), .en_x(wire_59[0:0]), .color_info(wire_69), .pixel_info(wire_59));
  TC_DotMatrixDisplay # (.UUID(64'd4046095411372047939 ^ UUID)) DotMatrixDisplay_503 (.clk(clk), .rst(rst), .en_y(wire_17[0:0]), .en_x(wire_59[0:0]), .color_info(wire_17), .pixel_info(wire_59));
  TC_DotMatrixDisplay # (.UUID(64'd4125954542330108464 ^ UUID)) DotMatrixDisplay_504 (.clk(clk), .rst(rst), .en_y(wire_20[0:0]), .en_x(wire_59[0:0]), .color_info(wire_20), .pixel_info(wire_59));
  TC_DotMatrixDisplay # (.UUID(64'd1830364245155235777 ^ UUID)) DotMatrixDisplay_505 (.clk(clk), .rst(rst), .en_y(wire_53[0:0]), .en_x(wire_30[0:0]), .color_info(wire_53), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd935797118162805439 ^ UUID)) DotMatrixDisplay_506 (.clk(clk), .rst(rst), .en_y(wire_66[0:0]), .en_x(wire_30[0:0]), .color_info(wire_66), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd3589916040253227553 ^ UUID)) DotMatrixDisplay_507 (.clk(clk), .rst(rst), .en_y(wire_105[0:0]), .en_x(wire_30[0:0]), .color_info(wire_105), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd433540754432702537 ^ UUID)) DotMatrixDisplay_508 (.clk(clk), .rst(rst), .en_y(wire_40[0:0]), .en_x(wire_30[0:0]), .color_info(wire_40), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd3645379267831978614 ^ UUID)) DotMatrixDisplay_509 (.clk(clk), .rst(rst), .en_y(wire_69[0:0]), .en_x(wire_30[0:0]), .color_info(wire_69), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd447614014945677748 ^ UUID)) DotMatrixDisplay_510 (.clk(clk), .rst(rst), .en_y(wire_17[0:0]), .en_x(wire_30[0:0]), .color_info(wire_17), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd3441989151667490927 ^ UUID)) DotMatrixDisplay_511 (.clk(clk), .rst(rst), .en_y(wire_20[0:0]), .en_x(wire_30[0:0]), .color_info(wire_20), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd1031401386565850890 ^ UUID)) DotMatrixDisplay_512 (.clk(clk), .rst(rst), .en_y(wire_53[0:0]), .en_x(wire_57[0:0]), .color_info(wire_53), .pixel_info(wire_57));
  TC_DotMatrixDisplay # (.UUID(64'd902548838630036546 ^ UUID)) DotMatrixDisplay_513 (.clk(clk), .rst(rst), .en_y(wire_66[0:0]), .en_x(wire_57[0:0]), .color_info(wire_66), .pixel_info(wire_57));
  TC_DotMatrixDisplay # (.UUID(64'd4178833354364662069 ^ UUID)) DotMatrixDisplay_514 (.clk(clk), .rst(rst), .en_y(wire_105[0:0]), .en_x(wire_57[0:0]), .color_info(wire_105), .pixel_info(wire_57));
  TC_DotMatrixDisplay # (.UUID(64'd4299503541740510209 ^ UUID)) DotMatrixDisplay_515 (.clk(clk), .rst(rst), .en_y(wire_40[0:0]), .en_x(wire_57[0:0]), .color_info(wire_40), .pixel_info(wire_57));
  TC_DotMatrixDisplay # (.UUID(64'd2917522327301819948 ^ UUID)) DotMatrixDisplay_516 (.clk(clk), .rst(rst), .en_y(wire_69[0:0]), .en_x(wire_57[0:0]), .color_info(wire_69), .pixel_info(wire_57));
  TC_DotMatrixDisplay # (.UUID(64'd3673936914473092842 ^ UUID)) DotMatrixDisplay_517 (.clk(clk), .rst(rst), .en_y(wire_17[0:0]), .en_x(wire_57[0:0]), .color_info(wire_17), .pixel_info(wire_57));
  TC_DotMatrixDisplay # (.UUID(64'd483335405037895454 ^ UUID)) DotMatrixDisplay_518 (.clk(clk), .rst(rst), .en_y(wire_20[0:0]), .en_x(wire_57[0:0]), .color_info(wire_20), .pixel_info(wire_57));
  TC_DotMatrixDisplay # (.UUID(64'd3207526772371322069 ^ UUID)) DotMatrixDisplay_519 (.clk(clk), .rst(rst), .en_y(wire_53[0:0]), .en_x(wire_33[0:0]), .color_info(wire_53), .pixel_info(wire_33));
  TC_DotMatrixDisplay # (.UUID(64'd856696257992628472 ^ UUID)) DotMatrixDisplay_520 (.clk(clk), .rst(rst), .en_y(wire_66[0:0]), .en_x(wire_33[0:0]), .color_info(wire_66), .pixel_info(wire_33));
  TC_DotMatrixDisplay # (.UUID(64'd1891245696899112287 ^ UUID)) DotMatrixDisplay_521 (.clk(clk), .rst(rst), .en_y(wire_105[0:0]), .en_x(wire_33[0:0]), .color_info(wire_105), .pixel_info(wire_33));
  TC_DotMatrixDisplay # (.UUID(64'd1832275632133913188 ^ UUID)) DotMatrixDisplay_522 (.clk(clk), .rst(rst), .en_y(wire_40[0:0]), .en_x(wire_33[0:0]), .color_info(wire_40), .pixel_info(wire_33));
  TC_DotMatrixDisplay # (.UUID(64'd2710136185812050848 ^ UUID)) DotMatrixDisplay_523 (.clk(clk), .rst(rst), .en_y(wire_69[0:0]), .en_x(wire_33[0:0]), .color_info(wire_69), .pixel_info(wire_33));
  TC_DotMatrixDisplay # (.UUID(64'd4572995742389431434 ^ UUID)) DotMatrixDisplay_524 (.clk(clk), .rst(rst), .en_y(wire_17[0:0]), .en_x(wire_33[0:0]), .color_info(wire_17), .pixel_info(wire_33));
  TC_DotMatrixDisplay # (.UUID(64'd1755821087589377818 ^ UUID)) DotMatrixDisplay_525 (.clk(clk), .rst(rst), .en_y(wire_20[0:0]), .en_x(wire_33[0:0]), .color_info(wire_20), .pixel_info(wire_33));
  TC_DotMatrixDisplay # (.UUID(64'd1516332879740996967 ^ UUID)) DotMatrixDisplay_526 (.clk(clk), .rst(rst), .en_y(wire_53[0:0]), .en_x(wire_2[0:0]), .color_info(wire_53), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd743797602559305145 ^ UUID)) DotMatrixDisplay_527 (.clk(clk), .rst(rst), .en_y(wire_66[0:0]), .en_x(wire_2[0:0]), .color_info(wire_66), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd1675081676777874763 ^ UUID)) DotMatrixDisplay_528 (.clk(clk), .rst(rst), .en_y(wire_105[0:0]), .en_x(wire_2[0:0]), .color_info(wire_105), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd1854067883140902272 ^ UUID)) DotMatrixDisplay_529 (.clk(clk), .rst(rst), .en_y(wire_40[0:0]), .en_x(wire_2[0:0]), .color_info(wire_40), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd4334581264551437851 ^ UUID)) DotMatrixDisplay_530 (.clk(clk), .rst(rst), .en_y(wire_69[0:0]), .en_x(wire_2[0:0]), .color_info(wire_69), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd1212294827969597911 ^ UUID)) DotMatrixDisplay_531 (.clk(clk), .rst(rst), .en_y(wire_17[0:0]), .en_x(wire_2[0:0]), .color_info(wire_17), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd4451864437363452741 ^ UUID)) DotMatrixDisplay_532 (.clk(clk), .rst(rst), .en_y(wire_20[0:0]), .en_x(wire_2[0:0]), .color_info(wire_20), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd660731318950632123 ^ UUID)) DotMatrixDisplay_533 (.clk(clk), .rst(rst), .en_y(wire_53[0:0]), .en_x(wire_47[0:0]), .color_info(wire_53), .pixel_info(wire_47));
  TC_DotMatrixDisplay # (.UUID(64'd3378460741643499424 ^ UUID)) DotMatrixDisplay_534 (.clk(clk), .rst(rst), .en_y(wire_66[0:0]), .en_x(wire_47[0:0]), .color_info(wire_66), .pixel_info(wire_47));
  TC_DotMatrixDisplay # (.UUID(64'd3603843643654745865 ^ UUID)) DotMatrixDisplay_535 (.clk(clk), .rst(rst), .en_y(wire_105[0:0]), .en_x(wire_47[0:0]), .color_info(wire_105), .pixel_info(wire_47));
  TC_DotMatrixDisplay # (.UUID(64'd2732406589031164731 ^ UUID)) DotMatrixDisplay_536 (.clk(clk), .rst(rst), .en_y(wire_40[0:0]), .en_x(wire_47[0:0]), .color_info(wire_40), .pixel_info(wire_47));
  TC_DotMatrixDisplay # (.UUID(64'd4137052652423786809 ^ UUID)) DotMatrixDisplay_537 (.clk(clk), .rst(rst), .en_y(wire_69[0:0]), .en_x(wire_47[0:0]), .color_info(wire_69), .pixel_info(wire_47));
  TC_DotMatrixDisplay # (.UUID(64'd1409126998886186295 ^ UUID)) DotMatrixDisplay_538 (.clk(clk), .rst(rst), .en_y(wire_17[0:0]), .en_x(wire_47[0:0]), .color_info(wire_17), .pixel_info(wire_47));
  TC_DotMatrixDisplay # (.UUID(64'd1577612092082569527 ^ UUID)) DotMatrixDisplay_539 (.clk(clk), .rst(rst), .en_y(wire_20[0:0]), .en_x(wire_47[0:0]), .color_info(wire_20), .pixel_info(wire_47));
  TC_DotMatrixDisplay # (.UUID(64'd1379213194016457817 ^ UUID)) DotMatrixDisplay_540 (.clk(clk), .rst(rst), .en_y(wire_53[0:0]), .en_x(wire_31[0:0]), .color_info(wire_53), .pixel_info(wire_31));
  TC_DotMatrixDisplay # (.UUID(64'd3741196406093988473 ^ UUID)) DotMatrixDisplay_541 (.clk(clk), .rst(rst), .en_y(wire_66[0:0]), .en_x(wire_31[0:0]), .color_info(wire_66), .pixel_info(wire_31));
  TC_DotMatrixDisplay # (.UUID(64'd2504220079177694680 ^ UUID)) DotMatrixDisplay_542 (.clk(clk), .rst(rst), .en_y(wire_105[0:0]), .en_x(wire_31[0:0]), .color_info(wire_105), .pixel_info(wire_31));
  TC_DotMatrixDisplay # (.UUID(64'd1788238612100923660 ^ UUID)) DotMatrixDisplay_543 (.clk(clk), .rst(rst), .en_y(wire_40[0:0]), .en_x(wire_31[0:0]), .color_info(wire_40), .pixel_info(wire_31));
  TC_DotMatrixDisplay # (.UUID(64'd348123188284652061 ^ UUID)) DotMatrixDisplay_544 (.clk(clk), .rst(rst), .en_y(wire_69[0:0]), .en_x(wire_31[0:0]), .color_info(wire_69), .pixel_info(wire_31));
  TC_DotMatrixDisplay # (.UUID(64'd297947842881024910 ^ UUID)) DotMatrixDisplay_545 (.clk(clk), .rst(rst), .en_y(wire_17[0:0]), .en_x(wire_31[0:0]), .color_info(wire_17), .pixel_info(wire_31));
  TC_DotMatrixDisplay # (.UUID(64'd3187027233044946476 ^ UUID)) DotMatrixDisplay_546 (.clk(clk), .rst(rst), .en_y(wire_20[0:0]), .en_x(wire_31[0:0]), .color_info(wire_20), .pixel_info(wire_31));
  TC_DotMatrixDisplay # (.UUID(64'd3974021049520770448 ^ UUID)) DotMatrixDisplay_547 (.clk(clk), .rst(rst), .en_y(wire_73[0:0]), .en_x(wire_38[0:0]), .color_info(wire_73), .pixel_info(wire_38));
  TC_DotMatrixDisplay # (.UUID(64'd3011377408596684094 ^ UUID)) DotMatrixDisplay_548 (.clk(clk), .rst(rst), .en_y(wire_73[0:0]), .en_x(wire_46[0:0]), .color_info(wire_73), .pixel_info(wire_46));
  TC_DotMatrixDisplay # (.UUID(64'd787806192135834626 ^ UUID)) DotMatrixDisplay_549 (.clk(clk), .rst(rst), .en_y(wire_73[0:0]), .en_x(wire_16[0:0]), .color_info(wire_73), .pixel_info(wire_16));
  TC_DotMatrixDisplay # (.UUID(64'd2982830508915352400 ^ UUID)) DotMatrixDisplay_550 (.clk(clk), .rst(rst), .en_y(wire_73[0:0]), .en_x(wire_11[0:0]), .color_info(wire_73), .pixel_info(wire_11));
  TC_DotMatrixDisplay # (.UUID(64'd2287184674519851503 ^ UUID)) DotMatrixDisplay_551 (.clk(clk), .rst(rst), .en_y(wire_73[0:0]), .en_x(wire_65[0:0]), .color_info(wire_73), .pixel_info(wire_65));
  TC_DotMatrixDisplay # (.UUID(64'd4015847227853570513 ^ UUID)) DotMatrixDisplay_552 (.clk(clk), .rst(rst), .en_y(wire_73[0:0]), .en_x(wire_7[0:0]), .color_info(wire_73), .pixel_info(wire_7));
  TC_DotMatrixDisplay # (.UUID(64'd4608460365758742729 ^ UUID)) DotMatrixDisplay_553 (.clk(clk), .rst(rst), .en_y(wire_73[0:0]), .en_x(wire_52[0:0]), .color_info(wire_73), .pixel_info(wire_52));
  TC_DotMatrixDisplay # (.UUID(64'd126678022832142258 ^ UUID)) DotMatrixDisplay_554 (.clk(clk), .rst(rst), .en_y(wire_73[0:0]), .en_x(wire_41[0:0]), .color_info(wire_73), .pixel_info(wire_41));
  TC_DotMatrixDisplay # (.UUID(64'd2875975831960078979 ^ UUID)) DotMatrixDisplay_555 (.clk(clk), .rst(rst), .en_y(wire_73[0:0]), .en_x(wire_59[0:0]), .color_info(wire_73), .pixel_info(wire_59));
  TC_DotMatrixDisplay # (.UUID(64'd4007631186959209700 ^ UUID)) DotMatrixDisplay_556 (.clk(clk), .rst(rst), .en_y(wire_73[0:0]), .en_x(wire_30[0:0]), .color_info(wire_73), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd960426467855939903 ^ UUID)) DotMatrixDisplay_557 (.clk(clk), .rst(rst), .en_y(wire_73[0:0]), .en_x(wire_57[0:0]), .color_info(wire_73), .pixel_info(wire_57));
  TC_DotMatrixDisplay # (.UUID(64'd3269721929079556361 ^ UUID)) DotMatrixDisplay_558 (.clk(clk), .rst(rst), .en_y(wire_73[0:0]), .en_x(wire_33[0:0]), .color_info(wire_73), .pixel_info(wire_33));
  TC_DotMatrixDisplay # (.UUID(64'd1719689023077837617 ^ UUID)) DotMatrixDisplay_559 (.clk(clk), .rst(rst), .en_y(wire_73[0:0]), .en_x(wire_2[0:0]), .color_info(wire_73), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd966749569609805529 ^ UUID)) DotMatrixDisplay_560 (.clk(clk), .rst(rst), .en_y(wire_73[0:0]), .en_x(wire_47[0:0]), .color_info(wire_73), .pixel_info(wire_47));
  TC_Decoder3 # (.UUID(64'd1761087297263831232 ^ UUID)) Decoder3_561 (.dis(wire_29), .sel0(wire_167), .sel1(wire_39), .sel2(wire_200), .out0(wire_405), .out1(wire_122), .out2(wire_246), .out3(wire_454), .out4(wire_414), .out5(wire_382), .out6(wire_247), .out7(wire_442));
  TC_Or # (.UUID(64'd2054144748014383948 ^ UUID), .BIT_WIDTH(64'd64)) Or64_562 (.in0(wire_208), .in1(wire_24), .out(wire_46));
  TC_Or # (.UUID(64'd699363347671241607 ^ UUID), .BIT_WIDTH(64'd64)) Or64_563 (.in0(wire_82), .in1({{56{1'b0}}, wire_308 }), .out(wire_208));
  TC_Or # (.UUID(64'd1724882088379321674 ^ UUID), .BIT_WIDTH(64'd64)) Or64_564 (.in0(wire_445), .in1(wire_24), .out(wire_16));
  TC_Or # (.UUID(64'd3048379343391964044 ^ UUID), .BIT_WIDTH(64'd64)) Or64_565 (.in0(wire_82), .in1({{56{1'b0}}, wire_403 }), .out(wire_445));
  TC_Or # (.UUID(64'd2856211505080343582 ^ UUID), .BIT_WIDTH(64'd64)) Or64_566 (.in0(wire_107), .in1(wire_24), .out(wire_11));
  TC_Or # (.UUID(64'd4267532593049086930 ^ UUID), .BIT_WIDTH(64'd64)) Or64_567 (.in0(wire_82), .in1({{56{1'b0}}, wire_409 }), .out(wire_107));
  TC_Or # (.UUID(64'd1141295085411161283 ^ UUID), .BIT_WIDTH(64'd64)) Or64_568 (.in0(wire_201), .in1(wire_24), .out(wire_65));
  TC_Or # (.UUID(64'd2957732111256797719 ^ UUID), .BIT_WIDTH(64'd64)) Or64_569 (.in0(wire_82), .in1({{56{1'b0}}, wire_120 }), .out(wire_201));
  TC_Or # (.UUID(64'd3075550721366977453 ^ UUID), .BIT_WIDTH(64'd64)) Or64_570 (.in0(wire_427), .in1(wire_24), .out(wire_7));
  TC_Or # (.UUID(64'd2213041841753283622 ^ UUID), .BIT_WIDTH(64'd64)) Or64_571 (.in0(wire_82), .in1({{56{1'b0}}, wire_319 }), .out(wire_427));
  TC_Or # (.UUID(64'd2863405907234665898 ^ UUID), .BIT_WIDTH(64'd64)) Or64_572 (.in0(wire_169), .in1(wire_24), .out(wire_52));
  TC_Or # (.UUID(64'd2507246242342996184 ^ UUID), .BIT_WIDTH(64'd64)) Or64_573 (.in0(wire_82), .in1({{56{1'b0}}, wire_153 }), .out(wire_169));
  TC_Or # (.UUID(64'd3603024006464314277 ^ UUID), .BIT_WIDTH(64'd64)) Or64_574 (.in0(wire_300), .in1(wire_24), .out(wire_41));
  TC_Or # (.UUID(64'd4385757953256632425 ^ UUID), .BIT_WIDTH(64'd64)) Or64_575 (.in0(wire_82), .in1({{63{1'b0}}, wire_28 }), .out(wire_300));
  TC_Or # (.UUID(64'd1819355801877563735 ^ UUID), .BIT_WIDTH(64'd64)) Or64_576 (.in0(wire_85), .in1(wire_24), .out(wire_59));
  TC_Or # (.UUID(64'd4533565317199406216 ^ UUID), .BIT_WIDTH(64'd64)) Or64_577 (.in0(wire_82), .in1({{63{1'b0}}, wire_210 }), .out(wire_85));
  TC_Or # (.UUID(64'd1223415715719310412 ^ UUID), .BIT_WIDTH(64'd64)) Or64_578 (.in0(wire_14), .in1(wire_24), .out(wire_30));
  TC_Or # (.UUID(64'd3751925248603012706 ^ UUID), .BIT_WIDTH(64'd64)) Or64_579 (.in0(wire_82), .in1({{63{1'b0}}, wire_112 }), .out(wire_14));
  TC_Or # (.UUID(64'd498599112880254247 ^ UUID), .BIT_WIDTH(64'd64)) Or64_580 (.in0(wire_243), .in1(wire_24), .out(wire_57));
  TC_Or # (.UUID(64'd4593450324580406305 ^ UUID), .BIT_WIDTH(64'd64)) Or64_581 (.in0(wire_82), .in1({{63{1'b0}}, wire_163 }), .out(wire_243));
  TC_Or # (.UUID(64'd3597486187217176065 ^ UUID), .BIT_WIDTH(64'd64)) Or64_582 (.in0(wire_232), .in1(wire_24), .out(wire_33));
  TC_Or # (.UUID(64'd3750411725135472848 ^ UUID), .BIT_WIDTH(64'd64)) Or64_583 (.in0(wire_82), .in1({{63{1'b0}}, wire_282 }), .out(wire_232));
  TC_Or # (.UUID(64'd1803132865256732472 ^ UUID), .BIT_WIDTH(64'd64)) Or64_584 (.in0(wire_335), .in1(wire_24), .out(wire_2));
  TC_Or # (.UUID(64'd3618716379687564923 ^ UUID), .BIT_WIDTH(64'd64)) Or64_585 (.in0(wire_82), .in1({{63{1'b0}}, wire_212 }), .out(wire_335));
  TC_Or # (.UUID(64'd250960130892132493 ^ UUID), .BIT_WIDTH(64'd64)) Or64_586 (.in0(wire_211), .in1(wire_24), .out(wire_47));
  TC_Or # (.UUID(64'd3915095558091040469 ^ UUID), .BIT_WIDTH(64'd64)) Or64_587 (.in0(wire_82), .in1({{63{1'b0}}, wire_343 }), .out(wire_211));
  TC_Or # (.UUID(64'd3328487448535793322 ^ UUID), .BIT_WIDTH(64'd64)) Or64_588 (.in0(wire_257), .in1(wire_24), .out(wire_31));
  TC_Or # (.UUID(64'd474644107318055740 ^ UUID), .BIT_WIDTH(64'd64)) Or64_589 (.in0(wire_82), .in1({{63{1'b0}}, wire_362 }), .out(wire_257));
  TC_Decoder3 # (.UUID(64'd955964025727377334 ^ UUID)) Decoder3_590 (.dis(wire_466), .sel0(wire_167), .sel1(wire_39), .sel2(wire_200), .out0(wire_28), .out1(wire_210), .out2(wire_112), .out3(wire_163), .out4(wire_282), .out5(wire_212), .out6(wire_343), .out7(wire_362));
  TC_DotMatrixDisplay # (.UUID(64'd285004982822351210 ^ UUID)) DotMatrixDisplay_591 (.clk(clk), .rst(rst), .en_y(wire_111[0:0]), .en_x(wire_19[0:0]), .color_info(wire_111), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd4383693547521216392 ^ UUID)) DotMatrixDisplay_592 (.clk(clk), .rst(rst), .en_y(wire_6[0:0]), .en_x(wire_19[0:0]), .color_info(wire_6), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd2932794430774723144 ^ UUID)) DotMatrixDisplay_593 (.clk(clk), .rst(rst), .en_y(wire_67[0:0]), .en_x(wire_19[0:0]), .color_info(wire_67), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd3959184663079228471 ^ UUID)) DotMatrixDisplay_594 (.clk(clk), .rst(rst), .en_y(wire_44[0:0]), .en_x(wire_19[0:0]), .color_info(wire_44), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd3064203474842665995 ^ UUID)) DotMatrixDisplay_595 (.clk(clk), .rst(rst), .en_y(wire_49[0:0]), .en_x(wire_19[0:0]), .color_info(wire_49), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd2900133665642818493 ^ UUID)) DotMatrixDisplay_596 (.clk(clk), .rst(rst), .en_y(wire_71[0:0]), .en_x(wire_19[0:0]), .color_info(wire_71), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd2793684364763582065 ^ UUID)) DotMatrixDisplay_597 (.clk(clk), .rst(rst), .en_y(wire_1[0:0]), .en_x(wire_19[0:0]), .color_info(wire_1), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd571922125710398315 ^ UUID)) DotMatrixDisplay_598 (.clk(clk), .rst(rst), .en_y(wire_102[0:0]), .en_x(wire_19[0:0]), .color_info(wire_102), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd402893291715572801 ^ UUID)) DotMatrixDisplay_599 (.clk(clk), .rst(rst), .en_y(wire_113[0:0]), .en_x(wire_19[0:0]), .color_info(wire_113), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd1792536061057532060 ^ UUID)) DotMatrixDisplay_600 (.clk(clk), .rst(rst), .en_y(wire_42[0:0]), .en_x(wire_19[0:0]), .color_info(wire_42), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd2938658035630064687 ^ UUID)) DotMatrixDisplay_601 (.clk(clk), .rst(rst), .en_y(wire_13[0:0]), .en_x(wire_19[0:0]), .color_info(wire_13), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd3609446542549819354 ^ UUID)) DotMatrixDisplay_602 (.clk(clk), .rst(rst), .en_y(wire_92[0:0]), .en_x(wire_19[0:0]), .color_info(wire_92), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd1767128864166779932 ^ UUID)) DotMatrixDisplay_603 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_19[0:0]), .color_info(wire_22), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd2404036166266630994 ^ UUID)) DotMatrixDisplay_604 (.clk(clk), .rst(rst), .en_y(wire_45[0:0]), .en_x(wire_19[0:0]), .color_info(wire_45), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd2628550272356333812 ^ UUID)) DotMatrixDisplay_605 (.clk(clk), .rst(rst), .en_y(wire_53[0:0]), .en_x(wire_19[0:0]), .color_info(wire_53), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd2517404727507393468 ^ UUID)) DotMatrixDisplay_606 (.clk(clk), .rst(rst), .en_y(wire_66[0:0]), .en_x(wire_19[0:0]), .color_info(wire_66), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd189626427841181534 ^ UUID)) DotMatrixDisplay_607 (.clk(clk), .rst(rst), .en_y(wire_105[0:0]), .en_x(wire_19[0:0]), .color_info(wire_105), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd2973156979347166644 ^ UUID)) DotMatrixDisplay_608 (.clk(clk), .rst(rst), .en_y(wire_40[0:0]), .en_x(wire_19[0:0]), .color_info(wire_40), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd3387033223438399684 ^ UUID)) DotMatrixDisplay_609 (.clk(clk), .rst(rst), .en_y(wire_69[0:0]), .en_x(wire_19[0:0]), .color_info(wire_69), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd4317828538525984487 ^ UUID)) DotMatrixDisplay_610 (.clk(clk), .rst(rst), .en_y(wire_17[0:0]), .en_x(wire_19[0:0]), .color_info(wire_17), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd2546702078073420598 ^ UUID)) DotMatrixDisplay_611 (.clk(clk), .rst(rst), .en_y(wire_20[0:0]), .en_x(wire_19[0:0]), .color_info(wire_20), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd4578656265108279561 ^ UUID)) DotMatrixDisplay_612 (.clk(clk), .rst(rst), .en_y(wire_73[0:0]), .en_x(wire_19[0:0]), .color_info(wire_73), .pixel_info(wire_19));
  TC_Or # (.UUID(64'd1151169897315353566 ^ UUID), .BIT_WIDTH(64'd64)) Or64_613 (.in0(wire_109), .in1(wire_24), .out(wire_19));
  TC_Or # (.UUID(64'd3456062963413460022 ^ UUID), .BIT_WIDTH(64'd64)) Or64_614 (.in0({{56{1'b0}}, wire_459 }), .in1(wire_82), .out(wire_109));
  TC_Or # (.UUID(64'd1502826367580921037 ^ UUID), .BIT_WIDTH(64'd64)) Or64_615 (.in0(wire_82), .in1({{56{1'b0}}, wire_457 }), .out(wire_281));
  TC_Or # (.UUID(64'd1854759391724557696 ^ UUID), .BIT_WIDTH(64'd64)) Or64_616 (.in0(wire_24), .in1(wire_281), .out(wire_38));
  TC_Constant # (.UUID(64'd1258114333586888636 ^ UUID), .BIT_WIDTH(64'd64), .value(64'h100000000000000)) Constant64_617 (.out(wire_24));
  TC_DotMatrixDisplay # (.UUID(64'd3403094820525018166 ^ UUID)) DotMatrixDisplay_618 (.clk(clk), .rst(rst), .en_y(wire_111[0:0]), .en_x(wire_31[0:0]), .color_info(wire_111), .pixel_info(wire_31));
  TC_Or # (.UUID(64'd1480142637011528932 ^ UUID), .BIT_WIDTH(64'd32)) Or32_619 (.in0({{31{1'b0}}, wire_351 }), .in1(wire_3), .out(wire_111));
  TC_Or # (.UUID(64'd3283593169104501706 ^ UUID), .BIT_WIDTH(64'd32)) Or32_620 (.in0({{31{1'b0}}, wire_121 }), .in1(wire_3), .out(wire_6));
  TC_Or # (.UUID(64'd456310048193130579 ^ UUID), .BIT_WIDTH(64'd32)) Or32_621 (.in0({{31{1'b0}}, wire_422 }), .in1(wire_3), .out(wire_67));
  TC_Or # (.UUID(64'd954913857421913189 ^ UUID), .BIT_WIDTH(64'd32)) Or32_622 (.in0({{31{1'b0}}, wire_263 }), .in1(wire_3), .out(wire_44));
  TC_Or # (.UUID(64'd2053537699156809302 ^ UUID), .BIT_WIDTH(64'd32)) Or32_623 (.in0({{31{1'b0}}, wire_313 }), .in1(wire_3), .out(wire_49));
  TC_Or # (.UUID(64'd2293510296467188789 ^ UUID), .BIT_WIDTH(64'd32)) Or32_624 (.in0({{31{1'b0}}, wire_355 }), .in1(wire_3), .out(wire_71));
  TC_Or # (.UUID(64'd2687654398995872368 ^ UUID), .BIT_WIDTH(64'd32)) Or32_625 (.in0({{31{1'b0}}, wire_309 }), .in1(wire_3), .out(wire_1));
  TC_Or # (.UUID(64'd1348834436038662226 ^ UUID), .BIT_WIDTH(64'd32)) Or32_626 (.in0({{31{1'b0}}, wire_231 }), .in1(wire_3), .out(wire_102));
  TC_Or # (.UUID(64'd624204125600545237 ^ UUID), .BIT_WIDTH(64'd32)) Or32_627 (.in0({{31{1'b0}}, wire_393 }), .in1(wire_3), .out(wire_113));
  TC_Or # (.UUID(64'd3727009402301135636 ^ UUID), .BIT_WIDTH(64'd32)) Or32_628 (.in0({{31{1'b0}}, wire_174 }), .in1(wire_3), .out(wire_42));
  TC_Or # (.UUID(64'd335105193488601816 ^ UUID), .BIT_WIDTH(64'd32)) Or32_629 (.in0({{31{1'b0}}, wire_84 }), .in1(wire_3), .out(wire_13));
  TC_Or # (.UUID(64'd359636882149561109 ^ UUID), .BIT_WIDTH(64'd32)) Or32_630 (.in0({{31{1'b0}}, wire_358 }), .in1(wire_3), .out(wire_92));
  TC_Or # (.UUID(64'd290638062856828299 ^ UUID), .BIT_WIDTH(64'd32)) Or32_631 (.in0({{31{1'b0}}, wire_23 }), .in1(wire_3), .out(wire_22));
  TC_Or # (.UUID(64'd1077905158186754969 ^ UUID), .BIT_WIDTH(64'd32)) Or32_632 (.in0({{31{1'b0}}, wire_271 }), .in1(wire_3), .out(wire_45));
  TC_Or # (.UUID(64'd1957959648479470428 ^ UUID), .BIT_WIDTH(64'd32)) Or32_633 (.in0({{31{1'b0}}, wire_340 }), .in1(wire_3), .out(wire_53));
  TC_Or # (.UUID(64'd1184563183654810013 ^ UUID), .BIT_WIDTH(64'd32)) Or32_634 (.in0({{31{1'b0}}, wire_276 }), .in1(wire_3), .out(wire_66));
  TC_Or # (.UUID(64'd3425410741172848698 ^ UUID), .BIT_WIDTH(64'd32)) Or32_635 (.in0({{31{1'b0}}, wire_447 }), .in1(wire_3), .out(wire_105));
  TC_Or # (.UUID(64'd483802579628661529 ^ UUID), .BIT_WIDTH(64'd32)) Or32_636 (.in0({{31{1'b0}}, wire_216 }), .in1(wire_3), .out(wire_40));
  TC_Or # (.UUID(64'd597169164633599749 ^ UUID), .BIT_WIDTH(64'd32)) Or32_637 (.in0({{31{1'b0}}, wire_185 }), .in1(wire_3), .out(wire_69));
  TC_Or # (.UUID(64'd4333979782052380663 ^ UUID), .BIT_WIDTH(64'd32)) Or32_638 (.in0({{31{1'b0}}, wire_262 }), .in1(wire_3), .out(wire_17));
  TC_Or # (.UUID(64'd2911657004411041778 ^ UUID), .BIT_WIDTH(64'd32)) Or32_639 (.in0({{31{1'b0}}, wire_119 }), .in1(wire_3), .out(wire_20));
  TC_Or # (.UUID(64'd160714023732906080 ^ UUID), .BIT_WIDTH(64'd32)) Or32_640 (.in0({{31{1'b0}}, wire_306 }), .in1(wire_3), .out(wire_73));
  TC_Splitter16 # (.UUID(64'd2962161457275136525 ^ UUID)) Splitter16_641 (.in(16'd0), .out0(wire_61), .out1(wire_126));
  TC_Maker16 # (.UUID(64'd605457519861865191 ^ UUID)) Maker16_642 (.in0(wire_61), .in1(wire_126), .out(wire_428));
  TC_And # (.UUID(64'd346554494124357010 ^ UUID), .BIT_WIDTH(64'd8)) And8_643 (.in0(wire_61), .in1(wire_250), .out(wire_171));
  TC_Constant # (.UUID(64'd726334783467739359 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1F)) Constant8_644 (.out(wire_250));
  TC_Shr # (.UUID(64'd2681097512250917063 ^ UUID), .BIT_WIDTH(64'd16)) Shr16_645 (.in(wire_428), .shift(wire_368), .out(wire_230));
  TC_Mul # (.UUID(64'd2874338680899878686 ^ UUID), .BIT_WIDTH(64'd8)) DivMod8_646 (.in0(wire_230[7:0]), .in1(wire_369), .out0(wire_223), .out1(wire_0));
  TC_And # (.UUID(64'd1236180052746557107 ^ UUID), .BIT_WIDTH(64'd8)) And8_647 (.in0(8'd0), .in1(wire_171), .out(wire_278));
  TC_Shr # (.UUID(64'd2761608549933656332 ^ UUID), .BIT_WIDTH(64'd8)) Shr8_648 (.in(wire_171), .shift(wire_62), .out(wire_497));
  TC_Mul # (.UUID(64'd2346430598743616706 ^ UUID), .BIT_WIDTH(64'd8)) Mul8_649 (.in0(wire_397), .in1(wire_0), .out0(wire_365), .out1());
  TC_Constant # (.UUID(64'd2089594524788636478 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h5)) Constant8_650 (.out(wire_368));
  TC_Constant # (.UUID(64'd4246998549797875356 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h8)) Constant8_651 (.out(wire_397));
  TC_Constant # (.UUID(64'd568064456355297963 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6)) Constant8_652 (.out(wire_369));
  TC_Maker16 # (.UUID(64'd4212127281314114567 ^ UUID)) Maker16_653 (.in0(wire_223), .in1(wire_497), .out());
  TC_Constant # (.UUID(64'd2372065517434057092 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h3)) Constant8_654 (.out(wire_62));
  TC_Splitter64 # (.UUID(64'd2786940585684961897 ^ UUID)) Splitter64_655 (.in(wire_143), .out0(wire_459), .out1(wire_457), .out2(wire_308), .out3(wire_403), .out4(wire_409), .out5(wire_120), .out6(wire_319), .out7(wire_153));
  TC_Maker64 # (.UUID(64'd3902992438838927717 ^ UUID)) Maker64_656 (.in0({{7{1'b0}}, wire_405 }), .in1({{7{1'b0}}, wire_122 }), .in2({{7{1'b0}}, wire_246 }), .in3({{7{1'b0}}, wire_454 }), .in4({{7{1'b0}}, wire_414 }), .in5({{7{1'b0}}, wire_382 }), .in6({{7{1'b0}}, wire_247 }), .in7({{7{1'b0}}, wire_442 }), .out(wire_143));
  TC_IndexerBit # (.UUID(64'd3321700142543428847 ^ UUID), .INDEX(64'd4)) IndexerBit_657 (.in({{63{1'b0}}, wire_70 }), .out(wire_429));
  TC_IndexerBit # (.UUID(64'd3547200117221810686 ^ UUID), .INDEX(64'd5)) IndexerBit_658 (.in({{63{1'b0}}, wire_70 }), .out());
  TC_IndexerBit # (.UUID(64'd3199140956936685004 ^ UUID), .INDEX(64'd1)) IndexerBit_659 (.in({{63{1'b0}}, wire_70 }), .out(wire_448));
  TC_IndexerBit # (.UUID(64'd4453486239931898957 ^ UUID), .INDEX(64'd0)) IndexerBit_660 (.in({{63{1'b0}}, wire_70 }), .out(wire_236));
  TC_IndexerBit # (.UUID(64'd793475158729231589 ^ UUID), .INDEX(64'd2)) IndexerBit_661 (.in({{63{1'b0}}, wire_70 }), .out(wire_337));
  TC_IndexerBit # (.UUID(64'd4137363779186351422 ^ UUID), .INDEX(64'd3)) IndexerBit_662 (.in({{63{1'b0}}, wire_70 }), .out(wire_391));
  TC_Maker64 # (.UUID(64'd455323208973641798 ^ UUID)) Maker64_663 (.in0(8'd0), .in1(wire_377[7:0]), .in2(wire_438[7:0]), .in3(wire_381[7:0]), .in4(wire_316[7:0]), .in5(wire_314[7:0]), .in6(wire_244[7:0]), .in7(8'd0), .out(wire_379));
  TC_Decoder3 # (.UUID(64'd3488486536041038265 ^ UUID)) Decoder3_664 (.dis(wire_186), .sel0(wire_391), .sel1(wire_429), .sel2(1'd0), .out0(wire_172), .out1(wire_180), .out2(wire_317), .out3(wire_130), .out4(wire_140), .out5(wire_331), .out6(), .out7());
  TC_Switch # (.UUID(64'd1208546562597426695 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_665 (.en(wire_331), .in({{56{1'b0}}, wire_147 }), .out(wire_244));
  TC_Switch # (.UUID(64'd1352249394905457759 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_666 (.en(wire_140), .in({{56{1'b0}}, wire_147 }), .out(wire_314));
  TC_Switch # (.UUID(64'd1967225638606888144 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_667 (.en(wire_130), .in({{56{1'b0}}, wire_147 }), .out(wire_316));
  TC_Switch # (.UUID(64'd4315271759461120500 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_668 (.en(wire_317), .in({{56{1'b0}}, wire_147 }), .out(wire_381));
  TC_Switch # (.UUID(64'd2206888624251500513 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_669 (.en(wire_180), .in({{56{1'b0}}, wire_147 }), .out(wire_438));
  TC_Switch # (.UUID(64'd1473709270489726686 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_670 (.en(wire_172), .in({{56{1'b0}}, wire_147 }), .out(wire_377));
  TC_Maker8 # (.UUID(64'd2980779663314168059 ^ UUID)) Maker8_671 (.in0(wire_64), .in1(wire_434), .in2(wire_460), .in3(wire_461), .in4(wire_277), .in5(wire_204), .in6(wire_469), .in7(wire_280), .out(wire_147));
  TC_Decoder3 # (.UUID(64'd2084405174033346046 ^ UUID)) Decoder3_672 (.dis(1'd0), .sel0(wire_236), .sel1(wire_448), .sel2(wire_337), .out0(wire_64), .out1(wire_434), .out2(wire_460), .out3(wire_461), .out4(wire_277), .out5(wire_204), .out6(wire_469), .out7(wire_280));
  TC_IndexerBit # (.UUID(64'd491317431227122727 ^ UUID), .INDEX(64'd2)) IndexerBit_673 (.in({{48{1'b0}}, wire_81 }), .out(wire_162));
  TC_IndexerBit # (.UUID(64'd1784556959547968077 ^ UUID), .INDEX(64'd1)) IndexerBit_674 (.in({{48{1'b0}}, wire_81 }), .out(wire_242));
  TC_IndexerBit # (.UUID(64'd3918991488535010924 ^ UUID), .INDEX(64'd0)) IndexerBit_675 (.in({{48{1'b0}}, wire_81 }), .out(wire_287));
  TC_Decoder3 # (.UUID(64'd3328016767844708558 ^ UUID)) Decoder3_676 (.dis(wire_496), .sel0(wire_287), .sel1(wire_242), .sel2(wire_162), .out0(wire_447), .out1(wire_216), .out2(wire_185), .out3(wire_262), .out4(wire_119), .out5(wire_306), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd94465637011135503 ^ UUID)) Decoder3_677 (.dis(wire_89), .sel0(wire_287), .sel1(wire_242), .sel2(wire_162), .out0(wire_393), .out1(wire_174), .out2(wire_84), .out3(wire_358), .out4(wire_23), .out5(wire_271), .out6(wire_340), .out7(wire_276));
  TC_Decoder3 # (.UUID(64'd4134532680229405618 ^ UUID)) Decoder3_678 (.dis(wire_375), .sel0(wire_287), .sel1(wire_242), .sel2(wire_162), .out0(wire_351), .out1(wire_121), .out2(wire_422), .out3(wire_263), .out4(wire_313), .out5(wire_355), .out6(wire_309), .out7(wire_231));
  TC_IndexerBit # (.UUID(64'd1791468559137273491 ^ UUID), .INDEX(64'd4)) IndexerBit_679 (.in({{56{1'b0}}, wire_170 }), .out(wire_97));
  TC_IndexerBit # (.UUID(64'd39658275061510058 ^ UUID), .INDEX(64'd5)) IndexerBit_680 (.in({{56{1'b0}}, wire_170 }), .out(wire_480));
  TC_IndexerBit # (.UUID(64'd892425656436566477 ^ UUID), .INDEX(64'd1)) IndexerBit_681 (.in({{56{1'b0}}, wire_170 }), .out(wire_117));
  TC_IndexerBit # (.UUID(64'd1773248366378408484 ^ UUID), .INDEX(64'd0)) IndexerBit_682 (.in({{56{1'b0}}, wire_170 }), .out(wire_224));
  TC_IndexerBit # (.UUID(64'd4486692224417328602 ^ UUID), .INDEX(64'd2)) IndexerBit_683 (.in({{56{1'b0}}, wire_170 }), .out(wire_148));
  TC_IndexerBit # (.UUID(64'd2599804714622620522 ^ UUID), .INDEX(64'd3)) IndexerBit_684 (.in({{56{1'b0}}, wire_170 }), .out(wire_376));
  TC_Maker64 # (.UUID(64'd3840288022000377902 ^ UUID)) Maker64_685 (.in0(8'd0), .in1(wire_361), .in2(wire_256), .in3(wire_87), .in4(wire_285), .in5(wire_118), .in6(wire_225), .in7(8'd0), .out(wire_82));
  TC_Decoder3 # (.UUID(64'd3726668915122675664 ^ UUID)) Decoder3_686 (.dis(wire_32), .sel0(wire_376), .sel1(wire_97), .sel2(wire_480), .out0(wire_213), .out1(wire_336), .out2(wire_324), .out3(wire_198), .out4(wire_54), .out5(wire_283), .out6(), .out7());
  TC_Maker8 # (.UUID(64'd1198523190652649461 ^ UUID)) Maker8_687 (.in0(wire_15), .in1(wire_330), .in2(wire_402), .in3(wire_388), .in4(wire_406), .in5(wire_446), .in6(wire_315), .in7(wire_275), .out(wire_248));
  TC_Decoder3 # (.UUID(64'd3560160864540717355 ^ UUID)) Decoder3_688 (.dis(1'd0), .sel0(wire_224), .sel1(wire_117), .sel2(wire_148), .out0(wire_15), .out1(wire_330), .out2(wire_402), .out3(wire_388), .out4(wire_406), .out5(wire_446), .out6(wire_315), .out7(wire_275));
  TC_IndexerBit # (.UUID(64'd1141394094657830628 ^ UUID), .INDEX(64'd2)) IndexerBit_689 (.in({{56{1'b0}}, wire_176 }), .out(wire_200));
  TC_IndexerBit # (.UUID(64'd696455848819800145 ^ UUID), .INDEX(64'd1)) IndexerBit_690 (.in({{56{1'b0}}, wire_176 }), .out(wire_39));
  TC_IndexerBit # (.UUID(64'd4432442853893919896 ^ UUID), .INDEX(64'd0)) IndexerBit_691 (.in({{56{1'b0}}, wire_176 }), .out(wire_167));
  TC_Not # (.UUID(64'd4158174356767112018 ^ UUID), .BIT_WIDTH(64'd1)) Not_692 (.in(wire_29), .out(wire_466));
  TC_IndexerBit # (.UUID(64'd828437776429867100 ^ UUID), .INDEX(64'd3)) IndexerBit_693 (.in({{56{1'b0}}, wire_399 }), .out(wire_29));
  TC_Switch # (.UUID(64'd1242485156338857011 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_694 (.en(wire_213), .in(wire_248), .out(wire_361));
  TC_Switch # (.UUID(64'd2401145753266180686 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_695 (.en(wire_336), .in(wire_248), .out(wire_256));
  TC_Switch # (.UUID(64'd170148487718755518 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_696 (.en(wire_324), .in(wire_248), .out(wire_87));
  TC_Switch # (.UUID(64'd4356842233532369827 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_697 (.en(wire_198), .in(wire_248), .out(wire_285));
  TC_Switch # (.UUID(64'd281934008546165059 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_698 (.en(wire_54), .in(wire_248), .out(wire_118));
  TC_Switch # (.UUID(64'd2607951404340506150 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_699 (.en(wire_283), .in(wire_248), .out(wire_225));
  TC_Constant # (.UUID(64'd698311943952732907 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_700 (.out(wire_443));
  TC_Shl # (.UUID(64'd3454443531074987460 ^ UUID), .BIT_WIDTH(64'd8)) Shl8_701 (.in(wire_498), .shift(wire_443), .out(wire_349));
  TC_Constant # (.UUID(64'd1719458208507105480 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hF8)) Constant8_702 (.out(wire_482));
  TC_Shr # (.UUID(64'd1493084800744544313 ^ UUID), .BIT_WIDTH(64'd16)) Shr16_703 (.in(wire_160), .shift(wire_452), .out(wire_470));
  TC_And # (.UUID(64'd2411815527054584759 ^ UUID), .BIT_WIDTH(64'd8)) And8_704 (.in0(wire_470[7:0]), .in1(wire_332), .out(wire_134));
  TC_Shl # (.UUID(64'd3715701029303627047 ^ UUID), .BIT_WIDTH(64'd8)) Shl8_705 (.in(wire_234), .shift(wire_411), .out(wire_292));
  TC_Constant # (.UUID(64'd2987513562534289054 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h3)) Constant8_706 (.out(wire_411));
  TC_Splitter16 # (.UUID(64'd3466091847196817273 ^ UUID)) Splitter16_707 (.in(wire_160), .out0(wire_234), .out1(wire_498));
  TC_And # (.UUID(64'd4373000637541561499 ^ UUID), .BIT_WIDTH(64'd8)) And8_708 (.in0(wire_349), .in1(wire_482), .out(wire_182));
  TC_Constant # (.UUID(64'd394376885650305340 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hF8)) Constant8_709 (.out(wire_332));
  TC_Constant # (.UUID(64'd4541308606545096170 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h2)) Constant8_710 (.out(wire_452));
  TC_Equal # (.UUID(64'd1733416920015184194 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_711 (.in0(wire_78), .in1(wire_404), .out(wire_154));
  TC_Switch # (.UUID(64'd2423614426668088778 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_712 (.en(wire_154), .in(wire_51), .out(wire_160));
  TC_Or # (.UUID(64'd4586758808239302393 ^ UUID), .BIT_WIDTH(64'd1)) Or_713 (.in0(wire_154), .in1(wire_367), .out(wire_128));
  TC_Mux # (.UUID(64'd2760656294824721895 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_714 (.sel(wire_367), .in0(wire_345), .in1(16'd0), .out(wire_274));
  TC_Register # (.UUID(64'd3241586208636038889 ^ UUID), .BIT_WIDTH(64'd16)) Register16_715 (.clk(clk), .rst(rst), .load(wire_222), .save(wire_128), .in(wire_274), .out(wire_150));
  TC_Add # (.UUID(64'd4017916402226097699 ^ UUID), .BIT_WIDTH(64'd16)) Add16_716 (.in0(wire_150), .in1({{8{1'b0}}, wire_133 }), .ci(1'd0), .out(wire_345), .co());
  TC_Constant # (.UUID(64'd2312984758713823189 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_717 (.out(wire_133));
  TC_Constant # (.UUID(64'd2551553762740893708 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h9)) Constant8_718 (.out(wire_404));
  TC_Equal # (.UUID(64'd1636136138147839671 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_719 (.in0(wire_135), .in1(wire_78), .out(wire_367));
  TC_Splitter16 # (.UUID(64'd2307928026015545361 ^ UUID)) Splitter16_720 (.in(wire_150), .out0(wire_321), .out1());
  TC_And # (.UUID(64'd615602252699701093 ^ UUID), .BIT_WIDTH(64'd8)) And8_721 (.in0(wire_129), .in1(wire_321), .out(wire_371));
  TC_Constant # (.UUID(64'd131938052894061522 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7F)) Constant8_722 (.out(wire_129));
  TC_Shr # (.UUID(64'd2050246496933416059 ^ UUID), .BIT_WIDTH(64'd16)) Shr16_723 (.in(wire_150), .shift(wire_189), .out(wire_384));
  TC_And # (.UUID(64'd481511477473248332 ^ UUID), .BIT_WIDTH(64'd8)) And8_724 (.in0(wire_360), .in1(wire_371), .out(wire_209));
  TC_Constant # (.UUID(64'd586021271185525686 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7)) Constant8_725 (.out(wire_360));
  TC_Mul # (.UUID(64'd1830091154931166947 ^ UUID), .BIT_WIDTH(64'd8)) DivMod8_726 (.in0(wire_384[7:0]), .in1(wire_354), .out0(wire_341), .out1(wire_462));
  TC_Shr # (.UUID(64'd2165163288895893939 ^ UUID), .BIT_WIDTH(64'd8)) Shr8_727 (.in(wire_371), .shift(wire_363), .out(wire_9));
  TC_Constant # (.UUID(64'd200810733702508651 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h3)) Constant8_728 (.out(wire_363));
  TC_Constant # (.UUID(64'd1630083914111217771 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7)) Constant8_729 (.out(wire_189));
  TC_Constant # (.UUID(64'd2652383470314897644 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6)) Constant8_730 (.out(wire_354));
  TC_Maker16 # (.UUID(64'd1681437785098422899 ^ UUID)) Maker16_731 (.in0(wire_341), .in1(wire_9), .out(wire_81));
  TC_Or # (.UUID(64'd3292255105432469957 ^ UUID), .BIT_WIDTH(64'd8)) Or8_732 (.in0(wire_328), .in1(wire_493), .out(wire_170));
  TC_DotMatrixDisplay # (.UUID(64'd3447635075793531404 ^ UUID)) DotMatrixDisplay_733 (.clk(clk), .rst(rst), .en_y(wire_102[0:0]), .en_x(wire_52[0:0]), .color_info(wire_102), .pixel_info(wire_52));
  TC_DotMatrixDisplay # (.UUID(64'd2357004856211857231 ^ UUID)) DotMatrixDisplay_734 (.clk(clk), .rst(rst), .en_y(wire_113[0:0]), .en_x(wire_52[0:0]), .color_info(wire_113), .pixel_info(wire_52));
  TC_DotMatrixDisplay # (.UUID(64'd4312010944155206568 ^ UUID)) DotMatrixDisplay_735 (.clk(clk), .rst(rst), .en_y(wire_102[0:0]), .en_x(wire_41[0:0]), .color_info(wire_102), .pixel_info(wire_41));
  TC_DotMatrixDisplay # (.UUID(64'd3431047806447067432 ^ UUID)) DotMatrixDisplay_736 (.clk(clk), .rst(rst), .en_y(wire_42[0:0]), .en_x(wire_52[0:0]), .color_info(wire_42), .pixel_info(wire_52));
  TC_DotMatrixDisplay # (.UUID(64'd4390021466414828942 ^ UUID)) DotMatrixDisplay_737 (.clk(clk), .rst(rst), .en_y(wire_113[0:0]), .en_x(wire_41[0:0]), .color_info(wire_113), .pixel_info(wire_41));
  TC_DotMatrixDisplay # (.UUID(64'd15653221926004127 ^ UUID)) DotMatrixDisplay_738 (.clk(clk), .rst(rst), .en_y(wire_42[0:0]), .en_x(wire_41[0:0]), .color_info(wire_42), .pixel_info(wire_41));
  TC_DotMatrixDisplay # (.UUID(64'd1014206133768206220 ^ UUID)) DotMatrixDisplay_739 (.clk(clk), .rst(rst), .en_y(wire_13[0:0]), .en_x(wire_52[0:0]), .color_info(wire_13), .pixel_info(wire_52));
  TC_DotMatrixDisplay # (.UUID(64'd2849325852045589 ^ UUID)) DotMatrixDisplay_740 (.clk(clk), .rst(rst), .en_y(wire_13[0:0]), .en_x(wire_41[0:0]), .color_info(wire_13), .pixel_info(wire_41));
  TC_DotMatrixDisplay # (.UUID(64'd314241367863885600 ^ UUID)) DotMatrixDisplay_741 (.clk(clk), .rst(rst), .en_y(wire_92[0:0]), .en_x(wire_41[0:0]), .color_info(wire_92), .pixel_info(wire_41));
  TC_Splitter16 # (.UUID(64'd3753172574692329186 ^ UUID)) Splitter16_742 (.in(wire_21[15:0]), .out0(), .out1(wire_78));
  TC_Constant # (.UUID(64'd2478682750138065728 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_743 (.out(wire_222));
  TC_Constant # (.UUID(64'd1856657540721794823 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h8)) Constant8_744 (.out(wire_135));
  TC_IndexerBit # (.UUID(64'd886570659050850114 ^ UUID), .INDEX(64'd7)) IndexerBit_745 (.in({{56{1'b0}}, wire_170 }), .out(wire_32));
  TC_Maker8 # (.UUID(64'd3468027941936484802 ^ UUID)) Maker8_746 (.in0(1'd0), .in1(1'd0), .in2(1'd0), .in3(1'd0), .in4(1'd0), .in5(1'd0), .in6(1'd0), .in7(wire_98), .out(wire_493));
  TC_Add # (.UUID(64'd4511269672692838297 ^ UUID), .BIT_WIDTH(64'd8)) Add8_747 (.in0(wire_209), .in1(wire_441), .ci(1'd0), .out(wire_328), .co());
  TC_Mul # (.UUID(64'd3054815539910482189 ^ UUID), .BIT_WIDTH(64'd8)) Mul8_748 (.in0(wire_489), .in1(wire_462), .out0(wire_441), .out1());
  TC_Constant # (.UUID(64'd3748427549873790510 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h8)) Constant8_749 (.out(wire_489));
  TC_Not # (.UUID(64'd556700617730582781 ^ UUID), .BIT_WIDTH(64'd1)) Not_750 (.in(wire_154), .out(wire_98));
  TC_IndexerByte # (.UUID(64'd200316289509724975 ^ UUID), .INDEX(64'd1)) IndexerByte_751 (.in({{48{1'b0}}, wire_81 }), .out(wire_176));
  TC_IndexerByte # (.UUID(64'd4536831201350273311 ^ UUID), .INDEX(64'd1)) IndexerByte_752 (.in({{48{1'b0}}, wire_81 }), .out(wire_399));
  TC_Maker32 # (.UUID(64'd282397218342167008 ^ UUID)) Maker32_753 (.in0(8'd0), .in1(wire_292), .in2(wire_134), .in3(wire_182), .out(wire_3));
  TC_Constant # (.UUID(64'd1106323522140457504 ^ UUID), .BIT_WIDTH(64'd16), .value(16'h21)) Constant16_754 (.out());
  TC_Decoder2 # (.UUID(64'd1231552903151527218 ^ UUID)) Decoder2_755 (.sel0(wire_270), .sel1(wire_494), .out0(wire_188), .out1(wire_279), .out2(wire_238), .out3());
  TC_IndexerBit # (.UUID(64'd2398859089020989329 ^ UUID), .INDEX(64'd4)) IndexerBit_756 (.in({{48{1'b0}}, wire_81 }), .out(wire_494));
  TC_IndexerBit # (.UUID(64'd3359636226302588737 ^ UUID), .INDEX(64'd3)) IndexerBit_757 (.in({{48{1'b0}}, wire_81 }), .out(wire_270));
  TC_Not # (.UUID(64'd2665383657229755682 ^ UUID), .BIT_WIDTH(64'd1)) Not_758 (.in(wire_188), .out(wire_375));
  TC_Not # (.UUID(64'd4154487238976036286 ^ UUID), .BIT_WIDTH(64'd1)) Not_759 (.in(wire_279), .out(wire_89));
  TC_Not # (.UUID(64'd1465380410737539706 ^ UUID), .BIT_WIDTH(64'd1)) Not_760 (.in(wire_238), .out(wire_496));
  TC_DotMatrixDisplay # (.UUID(64'd1161980261539595991 ^ UUID)) DotMatrixDisplay_761 (.clk(clk), .rst(rst), .en_y(wire_73[0:0]), .en_x(wire_31[0:0]), .color_info(wire_73), .pixel_info(wire_31));

  wire [7:0] wire_0;
  wire [31:0] wire_1;
  wire [63:0] wire_2;
  wire [31:0] wire_3;
  wire [15:0] wire_4;
  wire [0:0] wire_5;
  wire [31:0] wire_6;
  wire [63:0] wire_7;
  wire [15:0] wire_8;
  wire [7:0] wire_9;
  wire [15:0] wire_10;
  wire [63:0] wire_11;
  wire [15:0] wire_12;
  wire [15:0] wire_12_0;
  wire [15:0] wire_12_1;
  assign wire_12 = wire_12_0|wire_12_1;
  wire [31:0] wire_13;
  wire [63:0] wire_14;
  wire [0:0] wire_15;
  wire [63:0] wire_16;
  wire [31:0] wire_17;
  wire [0:0] wire_18;
  wire [63:0] wire_19;
  wire [31:0] wire_20;
  wire [63:0] wire_21;
  wire [31:0] wire_22;
  wire [0:0] wire_23;
  wire [63:0] wire_24;
  wire [15:0] wire_25;
  wire [0:0] wire_26;
  wire [7:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [63:0] wire_30;
  wire [63:0] wire_31;
  wire [0:0] wire_32;
  wire [63:0] wire_33;
  wire [0:0] wire_34;
  wire [7:0] wire_35;
  wire [63:0] wire_36;
  wire [15:0] wire_37;
  wire [63:0] wire_38;
  wire [0:0] wire_39;
  wire [31:0] wire_40;
  wire [63:0] wire_41;
  wire [31:0] wire_42;
  wire [0:0] wire_43;
  wire [31:0] wire_44;
  wire [31:0] wire_45;
  wire [63:0] wire_46;
  wire [63:0] wire_47;
  wire [31:0] wire_48;
  wire [31:0] wire_49;
  wire [15:0] wire_50;
  wire [15:0] wire_50_0;
  wire [15:0] wire_50_1;
  wire [15:0] wire_50_2;
  assign wire_50 = wire_50_0|wire_50_1|wire_50_2;
  wire [15:0] wire_51;
  wire [15:0] wire_51_0;
  wire [15:0] wire_51_1;
  assign wire_51 = wire_51_0|wire_51_1;
  wire [63:0] wire_52;
  wire [31:0] wire_53;
  wire [0:0] wire_54;
  wire [15:0] wire_55;
  wire [15:0] wire_56;
  wire [63:0] wire_57;
  wire [0:0] wire_58;
  wire [63:0] wire_59;
  wire [0:0] wire_60;
  wire [7:0] wire_61;
  wire [7:0] wire_62;
  wire [0:0] wire_63;
  wire [0:0] wire_64;
  wire [63:0] wire_65;
  wire [31:0] wire_66;
  wire [31:0] wire_67;
  wire [0:0] wire_68;
  wire [31:0] wire_69;
  wire [0:0] wire_70;
  assign wire_70 = 0;
  wire [31:0] wire_71;
  wire [0:0] wire_72;
  wire [31:0] wire_73;
  wire [15:0] wire_74;
  wire [0:0] wire_75;
  wire [15:0] wire_76;
  wire [0:0] wire_77;
  wire [7:0] wire_78;
  wire [15:0] wire_79;
  wire [15:0] wire_79_0;
  wire [15:0] wire_79_1;
  assign wire_79 = wire_79_0|wire_79_1;
  wire [15:0] wire_80;
  wire [15:0] wire_81;
  wire [63:0] wire_82;
  wire [63:0] wire_83;
  wire [63:0] wire_83_0;
  wire [63:0] wire_83_1;
  wire [63:0] wire_83_2;
  wire [63:0] wire_83_3;
  wire [63:0] wire_83_4;
  wire [63:0] wire_83_5;
  wire [63:0] wire_83_6;
  wire [63:0] wire_83_7;
  wire [63:0] wire_83_8;
  wire [63:0] wire_83_9;
  wire [63:0] wire_83_10;
  wire [63:0] wire_83_11;
  wire [63:0] wire_83_12;
  wire [63:0] wire_83_13;
  wire [63:0] wire_83_14;
  wire [63:0] wire_83_15;
  wire [63:0] wire_83_16;
  wire [63:0] wire_83_17;
  wire [63:0] wire_83_18;
  wire [63:0] wire_83_19;
  wire [63:0] wire_83_20;
  assign wire_83 = wire_83_0|wire_83_1|wire_83_2|wire_83_3|wire_83_4|wire_83_5|wire_83_6|wire_83_7|wire_83_8|wire_83_9|wire_83_10|wire_83_11|wire_83_12|wire_83_13|wire_83_14|wire_83_15|wire_83_16|wire_83_17|wire_83_18|wire_83_19|wire_83_20;
  wire [0:0] wire_84;
  wire [63:0] wire_85;
  wire [0:0] wire_86;
  wire [7:0] wire_87;
  wire [0:0] wire_88;
  wire [0:0] wire_89;
  wire [0:0] wire_90;
  wire [0:0] wire_90_0;
  wire [0:0] wire_90_1;
  wire [0:0] wire_90_2;
  wire [0:0] wire_90_3;
  wire [0:0] wire_90_4;
  wire [0:0] wire_90_5;
  wire [0:0] wire_90_6;
  wire [0:0] wire_90_7;
  wire [0:0] wire_90_8;
  wire [0:0] wire_90_9;
  assign wire_90 = wire_90_0|wire_90_1|wire_90_2|wire_90_3|wire_90_4|wire_90_5|wire_90_6|wire_90_7|wire_90_8|wire_90_9;
  wire [0:0] wire_91;
  wire [31:0] wire_92;
  wire [0:0] wire_93;
  wire [0:0] wire_94;
  wire [15:0] wire_95;
  wire [0:0] wire_96;
  wire [0:0] wire_97;
  wire [0:0] wire_98;
  wire [0:0] wire_99;
  wire [0:0] wire_100;
  wire [0:0] wire_100_0;
  wire [0:0] wire_100_1;
  wire [0:0] wire_100_2;
  assign wire_100 = wire_100_0|wire_100_1|wire_100_2;
  wire [15:0] wire_101;
  wire [31:0] wire_102;
  wire [7:0] wire_103;
  wire [63:0] wire_104;
  wire [31:0] wire_105;
  wire [15:0] wire_106;
  wire [63:0] wire_107;
  wire [7:0] wire_108;
  wire [63:0] wire_109;
  wire [0:0] wire_110;
  wire [31:0] wire_111;
  wire [0:0] wire_112;
  wire [31:0] wire_113;
  wire [0:0] wire_114;
  wire [0:0] wire_115;
  wire [7:0] wire_116;
  wire [0:0] wire_117;
  wire [7:0] wire_118;
  wire [0:0] wire_119;
  wire [7:0] wire_120;
  wire [0:0] wire_121;
  wire [0:0] wire_122;
  wire [15:0] wire_123;
  wire [0:0] wire_124;
  wire [0:0] wire_125;
  wire [7:0] wire_126;
  wire [0:0] wire_127;
  wire [0:0] wire_128;
  wire [7:0] wire_129;
  wire [0:0] wire_130;
  wire [0:0] wire_131;
  wire [0:0] wire_132;
  wire [7:0] wire_133;
  wire [7:0] wire_134;
  wire [7:0] wire_135;
  wire [15:0] wire_136;
  wire [0:0] wire_137;
  wire [0:0] wire_138;
  wire [0:0] wire_139;
  wire [0:0] wire_140;
  wire [0:0] wire_141;
  wire [0:0] wire_142;
  wire [63:0] wire_143;
  wire [0:0] wire_144;
  wire [0:0] wire_145;
  wire [0:0] wire_146;
  wire [7:0] wire_147;
  wire [0:0] wire_148;
  wire [15:0] wire_149;
  wire [15:0] wire_150;
  wire [15:0] wire_151;
  wire [0:0] wire_152;
  wire [7:0] wire_153;
  wire [0:0] wire_154;
  wire [15:0] wire_155;
  wire [0:0] wire_156;
  wire [0:0] wire_157;
  wire [0:0] wire_158;
  wire [0:0] wire_159;
  wire [15:0] wire_160;
  wire [0:0] wire_161;
  wire [0:0] wire_162;
  wire [0:0] wire_163;
  wire [7:0] wire_164;
  wire [0:0] wire_165;
  wire [0:0] wire_166;
  wire [0:0] wire_167;
  wire [15:0] wire_168;
  wire [63:0] wire_169;
  wire [7:0] wire_170;
  wire [7:0] wire_171;
  wire [0:0] wire_172;
  wire [15:0] wire_173;
  wire [0:0] wire_174;
  wire [0:0] wire_175;
  wire [7:0] wire_176;
  wire [15:0] wire_177;
  wire [0:0] wire_178;
  wire [15:0] wire_179;
  wire [0:0] wire_180;
  wire [0:0] wire_181;
  wire [7:0] wire_182;
  wire [0:0] wire_183;
  wire [15:0] wire_184;
  wire [0:0] wire_185;
  wire [0:0] wire_186;
  assign wire_186 = 0;
  wire [15:0] wire_187;
  wire [0:0] wire_188;
  wire [7:0] wire_189;
  wire [15:0] wire_190;
  wire [0:0] wire_191;
  wire [0:0] wire_192;
  wire [0:0] wire_193;
  wire [15:0] wire_194;
  wire [15:0] wire_194_0;
  wire [15:0] wire_194_1;
  assign wire_194 = wire_194_0|wire_194_1;
  wire [0:0] wire_195;
  wire [0:0] wire_196;
  wire [7:0] wire_197;
  wire [0:0] wire_198;
  wire [7:0] wire_199;
  wire [0:0] wire_200;
  wire [63:0] wire_201;
  wire [7:0] wire_202;
  wire [0:0] wire_203;
  wire [0:0] wire_204;
  wire [0:0] wire_205;
  wire [15:0] wire_206;
  wire [15:0] wire_207;
  wire [63:0] wire_208;
  wire [7:0] wire_209;
  wire [0:0] wire_210;
  wire [63:0] wire_211;
  wire [0:0] wire_212;
  wire [0:0] wire_213;
  wire [7:0] wire_214;
  wire [0:0] wire_215;
  wire [0:0] wire_216;
  wire [15:0] wire_217;
  wire [0:0] wire_218;
  wire [0:0] wire_219;
  wire [0:0] wire_220;
  wire [0:0] wire_221;
  wire [0:0] wire_222;
  wire [7:0] wire_223;
  wire [0:0] wire_224;
  wire [7:0] wire_225;
  wire [0:0] wire_226;
  wire [0:0] wire_227;
  wire [0:0] wire_228;
  wire [0:0] wire_229;
  wire [15:0] wire_230;
  wire [0:0] wire_231;
  wire [63:0] wire_232;
  wire [63:0] wire_233;
  wire [7:0] wire_234;
  wire [7:0] wire_235;
  wire [0:0] wire_236;
  wire [0:0] wire_237;
  wire [0:0] wire_238;
  wire [7:0] wire_239;
  wire [0:0] wire_240;
  wire [0:0] wire_241;
  wire [0:0] wire_242;
  wire [63:0] wire_243;
  wire [63:0] wire_244;
  wire [7:0] wire_245;
  wire [0:0] wire_246;
  wire [0:0] wire_247;
  wire [7:0] wire_248;
  wire [0:0] wire_249;
  wire [7:0] wire_250;
  wire [0:0] wire_251;
  wire [0:0] wire_252;
  wire [7:0] wire_253;
  wire [0:0] wire_254;
  wire [0:0] wire_255;
  wire [7:0] wire_256;
  wire [63:0] wire_257;
  wire [0:0] wire_258;
  wire [0:0] wire_259;
  wire [0:0] wire_260;
  wire [0:0] wire_261;
  wire [0:0] wire_262;
  wire [0:0] wire_263;
  wire [0:0] wire_264;
  wire [0:0] wire_265;
  wire [0:0] wire_266;
  wire [0:0] wire_267;
  wire [0:0] wire_268;
  wire [7:0] wire_269;
  wire [0:0] wire_270;
  wire [0:0] wire_271;
  wire [7:0] wire_272;
  wire [7:0] wire_273;
  wire [15:0] wire_274;
  wire [0:0] wire_275;
  wire [0:0] wire_276;
  wire [0:0] wire_277;
  wire [7:0] wire_278;
  wire [0:0] wire_279;
  wire [0:0] wire_280;
  wire [63:0] wire_281;
  wire [0:0] wire_282;
  wire [0:0] wire_283;
  wire [0:0] wire_284;
  wire [7:0] wire_285;
  wire [0:0] wire_286;
  wire [0:0] wire_287;
  wire [15:0] wire_288;
  wire [15:0] wire_289;
  wire [15:0] wire_290;
  wire [0:0] wire_291;
  wire [7:0] wire_292;
  wire [15:0] wire_293;
  wire [63:0] wire_294;
  wire [0:0] wire_295;
  wire [0:0] wire_296;
  wire [0:0] wire_297;
  wire [15:0] wire_298;
  wire [0:0] wire_299;
  wire [63:0] wire_300;
  wire [0:0] wire_301;
  wire [0:0] wire_302;
  wire [15:0] wire_303;
  wire [0:0] wire_304;
  wire [0:0] wire_305;
  wire [0:0] wire_306;
  wire [0:0] wire_307;
  wire [7:0] wire_308;
  wire [0:0] wire_309;
  wire [0:0] wire_310;
  wire [15:0] wire_311;
  wire [15:0] wire_312;
  wire [0:0] wire_313;
  wire [63:0] wire_314;
  wire [0:0] wire_315;
  wire [63:0] wire_316;
  wire [0:0] wire_317;
  wire [0:0] wire_318;
  wire [7:0] wire_319;
  wire [7:0] wire_320;
  wire [7:0] wire_321;
  wire [0:0] wire_322;
  wire [0:0] wire_323;
  wire [0:0] wire_324;
  wire [0:0] wire_325;
  wire [15:0] wire_326;
  wire [63:0] wire_327;
  wire [7:0] wire_328;
  wire [0:0] wire_329;
  wire [0:0] wire_330;
  wire [0:0] wire_331;
  wire [7:0] wire_332;
  wire [0:0] wire_333;
  wire [0:0] wire_334;
  wire [63:0] wire_335;
  wire [0:0] wire_336;
  wire [0:0] wire_337;
  wire [0:0] wire_338;
  assign arch_output_enable = wire_338;
  wire [0:0] wire_339;
  wire [0:0] wire_340;
  wire [7:0] wire_341;
  wire [0:0] wire_342;
  wire [0:0] wire_343;
  wire [7:0] wire_344;
  wire [15:0] wire_345;
  wire [15:0] wire_346;
  wire [0:0] wire_347;
  wire [15:0] wire_348;
  wire [7:0] wire_349;
  wire [0:0] wire_350;
  wire [0:0] wire_351;
  wire [0:0] wire_352;
  wire [15:0] wire_353;
  wire [7:0] wire_354;
  wire [0:0] wire_355;
  wire [0:0] wire_356;
  wire [0:0] wire_357;
  wire [0:0] wire_358;
  wire [63:0] wire_359;
  wire [7:0] wire_360;
  wire [7:0] wire_361;
  wire [0:0] wire_362;
  wire [7:0] wire_363;
  wire [7:0] wire_364;
  wire [7:0] wire_365;
  wire [15:0] wire_366;
  wire [0:0] wire_367;
  wire [7:0] wire_368;
  wire [7:0] wire_369;
  wire [0:0] wire_370;
  wire [7:0] wire_371;
  wire [0:0] wire_372;
  wire [0:0] wire_373;
  wire [0:0] wire_374;
  wire [0:0] wire_375;
  wire [0:0] wire_376;
  wire [63:0] wire_377;
  wire [0:0] wire_378;
  wire [63:0] wire_379;
  wire [15:0] wire_380;
  wire [63:0] wire_381;
  wire [0:0] wire_382;
  wire [0:0] wire_383;
  wire [15:0] wire_384;
  wire [7:0] wire_385;
  wire [0:0] wire_386;
  wire [0:0] wire_387;
  wire [0:0] wire_388;
  wire [15:0] wire_389;
  wire [15:0] wire_390;
  wire [0:0] wire_391;
  wire [15:0] wire_392;
  wire [0:0] wire_393;
  wire [0:0] wire_394;
  assign wire_394 = 0;
  wire [15:0] wire_395;
  wire [0:0] wire_396;
  wire [7:0] wire_397;
  wire [0:0] wire_398;
  assign arch_input_enable = wire_398;
  wire [7:0] wire_399;
  wire [0:0] wire_400;
  wire [15:0] wire_401;
  wire [0:0] wire_402;
  wire [7:0] wire_403;
  wire [7:0] wire_404;
  wire [0:0] wire_405;
  wire [0:0] wire_406;
  wire [0:0] wire_407;
  wire [0:0] wire_408;
  wire [7:0] wire_409;
  wire [0:0] wire_410;
  wire [7:0] wire_411;
  wire [15:0] wire_412;
  wire [0:0] wire_413;
  wire [0:0] wire_414;
  wire [0:0] wire_415;
  wire [7:0] wire_416;
  wire [0:0] wire_417;
  wire [0:0] wire_418;
  wire [7:0] wire_419;
  wire [0:0] wire_420;
  wire [15:0] wire_421;
  wire [0:0] wire_422;
  wire [0:0] wire_423;
  wire [63:0] wire_424;
  wire [7:0] wire_425;
  wire [0:0] wire_426;
  wire [63:0] wire_427;
  wire [15:0] wire_428;
  wire [0:0] wire_429;
  wire [0:0] wire_430;
  wire [7:0] wire_431;
  wire [0:0] wire_432;
  wire [0:0] wire_433;
  wire [0:0] wire_434;
  wire [0:0] wire_435;
  wire [7:0] wire_436;
  wire [7:0] wire_437;
  wire [63:0] wire_438;
  wire [15:0] wire_439;
  wire [0:0] wire_440;
  wire [7:0] wire_441;
  wire [0:0] wire_442;
  wire [7:0] wire_443;
  wire [7:0] wire_444;
  wire [63:0] wire_445;
  wire [0:0] wire_446;
  wire [0:0] wire_447;
  wire [0:0] wire_448;
  wire [0:0] wire_449;
  wire [7:0] wire_450;
  wire [0:0] wire_451;
  wire [7:0] wire_452;
  wire [0:0] wire_453;
  wire [0:0] wire_454;
  wire [0:0] wire_455;
  wire [0:0] wire_456;
  wire [7:0] wire_457;
  wire [7:0] wire_458;
  wire [7:0] wire_459;
  wire [0:0] wire_460;
  wire [0:0] wire_461;
  wire [7:0] wire_462;
  wire [0:0] wire_463;
  wire [0:0] wire_464;
  wire [0:0] wire_465;
  wire [0:0] wire_466;
  wire [7:0] wire_467;
  wire [0:0] wire_468;
  wire [0:0] wire_469;
  wire [15:0] wire_470;
  wire [7:0] wire_471;
  wire [7:0] wire_472;
  wire [0:0] wire_473;
  wire [63:0] wire_474;
  wire [0:0] wire_475;
  wire [7:0] wire_476;
  wire [15:0] wire_477;
  wire [0:0] wire_478;
  wire [0:0] wire_479;
  wire [0:0] wire_480;
  wire [0:0] wire_481;
  wire [7:0] wire_482;
  wire [7:0] wire_483;
  wire [7:0] wire_484;
  wire [0:0] wire_485;
  wire [15:0] wire_486;
  wire [7:0] wire_487;
  wire [15:0] wire_488;
  wire [7:0] wire_489;
  wire [15:0] wire_490;
  wire [63:0] wire_491;
  wire [0:0] wire_492;
  wire [7:0] wire_493;
  wire [0:0] wire_494;
  wire [0:0] wire_495;
  wire [0:0] wire_496;
  wire [7:0] wire_497;
  wire [7:0] wire_498;

endmodule
