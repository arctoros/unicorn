module Unicornz_32x32 (clk, rst, arch_output_enable, arch_output_value, arch_input_enable, arch_input_value);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  output  wire [0:0] arch_output_enable;
  output  wire [7:0] arch_output_value;
  output  wire [0:0] arch_input_enable;
  input  wire [7:0] arch_input_value;

  TC_Program # (.UUID(64'd2054094413772625173 ^ UUID), .WORD_WIDTH(64'd16), .DEFAULT_FILE_NAME("Program_1C819BFC7C081515.w16.bin"), .ARG_SIG("Program_1C819BFC7C081515=%s")) Program_0 (.clk(clk), .rst(rst), .address(wire_312), .out0(wire_10), .out1(wire_126), .out2(wire_153), .out3(wire_143));
  TC_Decoder3 # (.UUID(64'd2564548179517358600 ^ UUID)) Decoder3_1 (.dis(wire_120), .sel0(wire_14), .sel1(wire_99), .sel2(wire_25), .out0(wire_26), .out1(wire_194), .out2(wire_174), .out3(wire_363), .out4(wire_284), .out5(wire_133), .out6(wire_362), .out7(wire_246));
  TC_Decoder3 # (.UUID(64'd3856915764158948127 ^ UUID)) Decoder3_2 (.dis(wire_295), .sel0(wire_14), .sel1(wire_99), .sel2(wire_25), .out0(wire_389), .out1(wire_302), .out2(wire_326), .out3(wire_385), .out4(wire_266), .out5(wire_94), .out6(wire_80), .out7(wire_157));
  TC_Decoder3 # (.UUID(64'd469263968959042607 ^ UUID)) Decoder3_3 (.dis(wire_337), .sel0(wire_14), .sel1(wire_99), .sel2(wire_25), .out0(wire_261), .out1(wire_145), .out2(wire_344), .out3(wire_262), .out4(wire_288), .out5(wire_91), .out6(wire_350), .out7(wire_264));
  TC_Decoder3 # (.UUID(64'd2355515313084503399 ^ UUID)) Decoder3_4 (.dis(wire_232), .sel0(wire_14), .sel1(wire_99), .sel2(wire_25), .out0(wire_238), .out1(wire_317), .out2(wire_405), .out3(wire_353), .out4(wire_115), .out5(wire_315), .out6(wire_382), .out7(wire_377));
  TC_Maker8 # (.UUID(64'd3412742270897961611 ^ UUID)) Maker8_5 (.in0(wire_26), .in1(wire_194), .in2(wire_174), .in3(wire_363), .in4(wire_284), .in5(wire_133), .in6(wire_362), .in7(wire_246), .out(wire_96));
  TC_Maker8 # (.UUID(64'd2545466735680713447 ^ UUID)) Maker8_6 (.in0(wire_389), .in1(wire_302), .in2(wire_326), .in3(wire_385), .in4(wire_266), .in5(wire_94), .in6(wire_80), .in7(wire_157), .out(wire_41));
  TC_Maker8 # (.UUID(64'd2498328128700172685 ^ UUID)) Maker8_7 (.in0(wire_261), .in1(wire_145), .in2(wire_344), .in3(wire_262), .in4(wire_288), .in5(wire_91), .in6(wire_350), .in7(wire_264), .out(wire_323));
  TC_Maker8 # (.UUID(64'd3307623088924666213 ^ UUID)) Maker8_8 (.in0(wire_238), .in1(wire_317), .in2(wire_405), .in3(wire_353), .in4(wire_115), .in5(wire_315), .in6(wire_382), .in7(wire_377), .out(wire_233));
  TC_Maker32 # (.UUID(64'd3223173008764962790 ^ UUID)) Maker32_9 (.in0(wire_233), .in1(wire_323), .in2(wire_41), .in3(wire_96), .out(wire_139));
  TC_Switch # (.UUID(64'd1126631217811470669 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_10 (.en(wire_298), .in(wire_136), .out(wire_161));
  TC_Switch # (.UUID(64'd383016835864160285 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_11 (.en(wire_18), .in(wire_132), .out(wire_35_0));
  TC_Switch # (.UUID(64'd3140243124393805415 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_12 (.en(wire_311), .in(wire_167), .out(wire_263));
  TC_Switch # (.UUID(64'd1581886471977480656 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_13 (.en(wire_114), .in(wire_167), .out(wire_97_0));
  TC_Switch # (.UUID(64'd2241249704231886051 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_14 (.en(wire_163), .in(wire_153[15:0]), .out(wire_132));
  TC_Switch # (.UUID(64'd4100643114395522594 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_15 (.en(wire_357), .in(wire_126[15:0]), .out(wire_136_1));
  TC_Switch # (.UUID(64'd8725165111331077 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_16 (.en(wire_273), .in(wire_153[15:0]), .out(wire_136_2));
  TC_Switch # (.UUID(64'd3499335185666676498 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_17 (.en(wire_163), .in(wire_143[15:0]), .out(wire_136_0));
  TC_And3 # (.UUID(64'd2537048141319315915 ^ UUID), .BIT_WIDTH(64'd1)) And3_18 (.in0(wire_213), .in1(wire_21), .in2(wire_220), .out(wire_13));
  TC_Program # (.UUID(64'd388994960009383908 ^ UUID), .WORD_WIDTH(64'd32), .DEFAULT_FILE_NAME("Program_565FCDAEAC6CFE4.w32.bin"), .ARG_SIG("Program_565FCDAEAC6CFE4=%s")) Program_19 (.clk(clk), .rst(rst), .address({{8{1'b0}}, wire_129 }), .out0(wire_83), .out1(), .out2(), .out3());
  TC_Not # (.UUID(64'd2992010998666944854 ^ UUID), .BIT_WIDTH(64'd1)) Not_20 (.in(wire_87), .out(wire_380));
  TC_Switch # (.UUID(64'd92717477479612822 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_21 (.en(wire_257), .in(wire_117), .out(wire_3));
  TC_Counter # (.UUID(64'd388538542796967315 ^ UUID), .BIT_WIDTH(64'd16), .count(16'd1)) Counter16_22 (.clk(clk), .rst(rst), .save(wire_87), .in(wire_86), .out(wire_144));
  TC_Counter # (.UUID(64'd3159443906265585347 ^ UUID), .BIT_WIDTH(64'd16), .count(16'd1)) Counter16_23 (.clk(clk), .rst(rst), .save(wire_287), .in(wire_86), .out(wire_66));
  TC_DelayLine # (.UUID(64'd1367561201104940128 ^ UUID), .BIT_WIDTH(64'd16)) DelayLine16_24 (.clk(clk), .rst(rst), .in(wire_1[15:0]), .out(wire_117));
  TC_Switch # (.UUID(64'd4093327232412684622 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_25 (.en(wire_87), .in(wire_66), .out(wire_98_1));
  TC_Switch # (.UUID(64'd3521663283135285715 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_26 (.en(wire_380), .in(wire_144), .out(wire_98_0));
  TC_Mux # (.UUID(64'd3040671060942591441 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_27 (.sel(wire_257), .in0(wire_98), .in1(wire_3), .out(wire_312));
  TC_DelayLine # (.UUID(64'd1970975974056862148 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_28 (.clk(clk), .rst(rst), .in(wire_54), .out(wire_257));
  TC_DelayLine # (.UUID(64'd4083747472069111906 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_29 (.clk(clk), .rst(rst), .in(wire_87), .out(wire_287));
  TC_Not # (.UUID(64'd2703499132143664233 ^ UUID), .BIT_WIDTH(64'd1)) Not_30 (.in(wire_287), .out(wire_87));
  TC_Not # (.UUID(64'd668729040907233308 ^ UUID), .BIT_WIDTH(64'd1)) Not_31 (.in(wire_25), .out(wire_392));
  TC_Not # (.UUID(64'd1492999759409908823 ^ UUID), .BIT_WIDTH(64'd1)) Not_32 (.in(wire_14), .out(wire_333));
  TC_And3 # (.UUID(64'd3485287916682882951 ^ UUID), .BIT_WIDTH(64'd1)) And3_33 (.in0(wire_392), .in1(wire_99), .in2(wire_333), .out(wire_220));
  TC_Switch # (.UUID(64'd1180978168546894742 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_34 (.en(wire_13), .in(wire_13), .out(wire_214_0));
  TC_Switch # (.UUID(64'd3723419762929890741 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_35 (.en(wire_273), .in(wire_273), .out(wire_214_1));
  TC_Switch # (.UUID(64'd2050768528734077835 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_36 (.en(wire_163), .in(wire_163), .out(wire_214_2));
  TC_Switch # (.UUID(64'd3057161046631511266 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_37 (.en(wire_251), .in(wire_251), .out(wire_273));
  TC_Decoder2 # (.UUID(64'd3508168605160458460 ^ UUID)) Decoder2_38 (.sel0(wire_281), .sel1(wire_171), .out0(), .out1(), .out2(wire_345), .out3(wire_251));
  TC_Not # (.UUID(64'd1768466669334456870 ^ UUID), .BIT_WIDTH(64'd1)) Not_39 (.in(wire_13), .out(wire_209));
  TC_Not # (.UUID(64'd3282289532960715218 ^ UUID), .BIT_WIDTH(64'd1)) Not_40 (.in(wire_88), .out(wire_295));
  TC_Not # (.UUID(64'd1327891776776277559 ^ UUID), .BIT_WIDTH(64'd1)) Not_41 (.in(wire_331), .out(wire_337));
  TC_Not # (.UUID(64'd1982359815710823425 ^ UUID), .BIT_WIDTH(64'd1)) Not_42 (.in(wire_130), .out(wire_232));
  TC_Decoder2 # (.UUID(64'd2605064451303635720 ^ UUID)) Decoder2_43 (.sel0(wire_21), .sel1(wire_213), .out0(wire_130), .out1(wire_331), .out2(wire_88), .out3(wire_334));
  TC_Add # (.UUID(64'd3313543325696297390 ^ UUID), .BIT_WIDTH(64'd16)) Add16_44 (.in0(wire_312), .in1(wire_83[15:0]), .ci(1'd0), .out(wire_86), .co());
  TC_IndexerBit # (.UUID(64'd2196806765189308211 ^ UUID), .INDEX(64'd1)) IndexerBit_45 (.in(wire_83), .out(wire_171));
  TC_IndexerBit # (.UUID(64'd737839460036088508 ^ UUID), .INDEX(64'd0)) IndexerBit_46 (.in(wire_83), .out(wire_281));
  TC_IndexerBit # (.UUID(64'd2903462054980356400 ^ UUID), .INDEX(64'd2)) IndexerBit_47 (.in(wire_83), .out(wire_163));
  TC_Splitter8 # (.UUID(64'd3910511016620535394 ^ UUID)) Splitter8_48 (.in(wire_347), .out0(wire_44), .out1(wire_67), .out2(wire_77), .out3(wire_31), .out4(wire_60), .out5(wire_200), .out6(wire_53), .out7(wire_111));
  TC_IndexerByte # (.UUID(64'd2436263972142084427 ^ UUID), .INDEX(64'd1)) IndexerByte_49 (.in({{32{1'b0}}, wire_139 }), .out(wire_347));
  TC_Switch # (.UUID(64'd607808644696146469 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_50 (.en(wire_44), .in(wire_242), .out(wire_1_2[15:0]));
  TC_Switch # (.UUID(64'd2632353714035774615 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_51 (.en(wire_67), .in(wire_369), .out(wire_1_5[15:0]));
  TC_Switch # (.UUID(64'd2222450423847071001 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_52 (.en(wire_77), .in(wire_125), .out(wire_1_8[15:0]));
  TC_Switch # (.UUID(64'd3314256307520299439 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_53 (.en(wire_31), .in(wire_280), .out(wire_1_10[15:0]));
  TC_Switch # (.UUID(64'd2595134878720988598 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_54 (.en(wire_60), .in(wire_181), .out(wire_1_12[15:0]));
  TC_Switch # (.UUID(64'd1299382207876995858 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_55 (.en(wire_200), .in(wire_147), .out(wire_1_14[15:0]));
  TC_Switch # (.UUID(64'd1287692551111612372 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_56 (.en(wire_53), .in(wire_305), .out(wire_1_16[15:0]));
  TC_Switch # (.UUID(64'd1141911395405296382 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_57 (.en(wire_111), .in({{8{1'b0}}, wire_278 }), .out(wire_1_17[15:0]));
  TC_Not # (.UUID(64'd3575339823787626444 ^ UUID), .BIT_WIDTH(64'd8)) Not8_58 (.in(wire_97[7:0]), .out(wire_278));
  TC_Rol # (.UUID(64'd2078177537373562034 ^ UUID), .BIT_WIDTH(64'd16)) Rol16_59 (.in(wire_97), .shift(wire_35[7:0]), .out(wire_305));
  TC_Shl # (.UUID(64'd4491813690601887022 ^ UUID), .BIT_WIDTH(64'd16)) Shl16_60 (.in(wire_97), .shift(wire_35[7:0]), .out(wire_181));
  TC_Shr # (.UUID(64'd4199576277751456538 ^ UUID), .BIT_WIDTH(64'd16)) Shr16_61 (.in(wire_97), .shift(wire_35[7:0]), .out(wire_280));
  TC_Xor # (.UUID(64'd1780129286836567965 ^ UUID), .BIT_WIDTH(64'd16)) Xor16_62 (.in0(wire_97), .in1(wire_35), .out(wire_125));
  TC_Or # (.UUID(64'd3629729579801707084 ^ UUID), .BIT_WIDTH(64'd16)) Or16_63 (.in0(wire_97), .in1(wire_35), .out(wire_369));
  TC_And # (.UUID(64'd3161317497787028707 ^ UUID), .BIT_WIDTH(64'd16)) And16_64 (.in0(wire_97), .in1(wire_35), .out(wire_242));
  TC_And # (.UUID(64'd381639147620396883 ^ UUID), .BIT_WIDTH(64'd8)) And8_65 (.in0(wire_390), .in1(wire_10[7:0]), .out(wire_129));
  TC_Or3 # (.UUID(64'd3488800466009071346 ^ UUID), .BIT_WIDTH(64'd1)) Or3_66 (.in0(wire_4), .in1(wire_20), .in2(wire_29), .out(wire_154));
  TC_Or # (.UUID(64'd800125638954551844 ^ UUID), .BIT_WIDTH(64'd1)) Or_67 (.in0(wire_82), .in1(wire_20), .out(wire_339));
  TC_Neg # (.UUID(64'd3923101654540497550 ^ UUID), .BIT_WIDTH(64'd16)) Neg16_68 (.in(wire_62), .out(wire_203));
  TC_Mux # (.UUID(64'd4466247896286800046 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_69 (.sel(wire_329), .in0(wire_203), .in1(wire_62), .out(wire_387));
  TC_Mux # (.UUID(64'd4573628848997923160 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_70 (.sel(wire_38), .in0({{8{1'b0}}, wire_236 }), .in1(wire_35), .out(wire_269));
  TC_Ashr # (.UUID(64'd2002805807653529301 ^ UUID), .BIT_WIDTH(64'd16)) Ashr16_71 (.in(wire_97), .shift(wire_35[7:0]), .out(wire_403));
  TC_Neg # (.UUID(64'd1410727121580829106 ^ UUID), .BIT_WIDTH(64'd16)) Neg16_72 (.in(wire_97), .out(wire_190));
  TC_Mul # (.UUID(64'd409697540344457906 ^ UUID), .BIT_WIDTH(64'd16)) DivMod16_73 (.in0(wire_97), .in1(wire_269), .out0(wire_341), .out1());
  TC_Mul # (.UUID(64'd4230356226461292418 ^ UUID), .BIT_WIDTH(64'd16)) Mul16_74 (.in0(wire_35), .in1(wire_97), .out0(wire_282), .out1());
  TC_Add # (.UUID(64'd1348307715225101930 ^ UUID), .BIT_WIDTH(64'd16)) Add16_75 (.in0(wire_387), .in1(wire_97), .ci(1'd0), .out(wire_383), .co());
  TC_Switch # (.UUID(64'd3604076901724081385 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_76 (.en(wire_356), .in(wire_190), .out(wire_1_1[15:0]));
  TC_Switch # (.UUID(64'd4522803089722429170 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_77 (.en(wire_38), .in(wire_341), .out(wire_1_3[15:0]));
  TC_Switch # (.UUID(64'd202434256468217393 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_78 (.en(wire_195), .in(wire_282), .out(wire_1_6[15:0]));
  TC_Switch # (.UUID(64'd981527730647914060 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_79 (.en(wire_154), .in(wire_383), .out(wire_1_9[15:0]));
  TC_IndexerByte # (.UUID(64'd4236276122307665751 ^ UUID), .INDEX(64'd0)) IndexerByte_80 (.in({{32{1'b0}}, wire_139 }), .out(wire_158));
  TC_Splitter8 # (.UUID(64'd4515369816812696921 ^ UUID)) Splitter8_81 (.in(wire_158), .out0(wire_29), .out1(wire_20), .out2(wire_195), .out3(wire_38), .out4(wire_356), .out5(wire_135), .out6(wire_82), .out7(wire_95));
  TC_Or # (.UUID(64'd3775589699623562439 ^ UUID), .BIT_WIDTH(64'd1)) Or_82 (.in0(wire_135), .in1(wire_82), .out(wire_4));
  TC_Or # (.UUID(64'd119900405875326486 ^ UUID), .BIT_WIDTH(64'd1)) Or_83 (.in0(wire_49), .in1(wire_47), .out(wire_277));
  TC_Add # (.UUID(64'd2771599484257026352 ^ UUID), .BIT_WIDTH(64'd16)) Add16_84 (.in0(wire_185), .in1(wire_307), .ci(1'd0), .out(wire_283), .co());
  TC_Mux # (.UUID(64'd1916750704823682311 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_85 (.sel(wire_5), .in0(wire_149), .in1(wire_161), .out(wire_74));
  TC_Switch # (.UUID(64'd110187611622282684 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_86 (.en(wire_186), .in(wire_218[15:0]), .out(wire_35_1));
  TC_Or # (.UUID(64'd1550338206798762433 ^ UUID), .BIT_WIDTH(64'd1)) Or_87 (.in0(wire_156), .in1(wire_0), .out(wire_393));
  TC_Switch # (.UUID(64'd1104805846581678264 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_88 (.en(wire_393), .in(wire_379[15:0]), .out(wire_97_1));
  TC_Or # (.UUID(64'd1973201053711173902 ^ UUID), .BIT_WIDTH(64'd1)) Or_89 (.in0(wire_0), .in1(wire_351), .out(wire_338));
  TC_And # (.UUID(64'd373051892767174731 ^ UUID), .BIT_WIDTH(64'd1)) And_90 (.in0(wire_207), .in1(wire_156), .out(wire_351));
  TC_Mux # (.UUID(64'd2189639269723513602 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_91 (.sel(wire_207), .in0(wire_28), .in1(wire_86), .out(wire_361));
  TC_Or3 # (.UUID(64'd4386189682368290849 ^ UUID), .BIT_WIDTH(64'd1)) Or3_92 (.in0(wire_0), .in1(wire_227), .in2(wire_207), .out(wire_366));
  TC_Nor # (.UUID(64'd3810192346818398090 ^ UUID), .BIT_WIDTH(64'd1)) Nor_93 (.in0(wire_366), .in1(wire_40), .out(wire_327));
  TC_Mux # (.UUID(64'd4107077995071586514 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_94 (.sel(wire_327), .in0(wire_361), .in1(wire_1[15:0]), .out(wire_179));
  TC_Switch # (.UUID(64'd1346494715147404059 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_95 (.en(wire_215), .in(wire_70), .out(wire_54_7));
  TC_Splitter8 # (.UUID(64'd3709071160935573773 ^ UUID)) Splitter8_96 (.in(wire_373), .out0(wire_192), .out1(wire_199), .out2(wire_51), .out3(wire_79), .out4(wire_378), .out5(wire_162), .out6(wire_215), .out7(wire_76));
  TC_Switch # (.UUID(64'd4272543595848591881 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_97 (.en(wire_199), .in(wire_299), .out(wire_54_0));
  TC_Switch # (.UUID(64'd2673250751246411725 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_98 (.en(wire_51), .in(wire_107), .out(wire_54_1));
  TC_Switch # (.UUID(64'd4158444071236719644 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_99 (.en(wire_79), .in(wire_243), .out(wire_54_3));
  TC_Switch # (.UUID(64'd1076960299062071464 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_100 (.en(wire_378), .in(wire_197), .out(wire_54_4));
  TC_Switch # (.UUID(64'd2871129963461955678 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_101 (.en(wire_162), .in(wire_206), .out(wire_54_6));
  TC_Switch # (.UUID(64'd1466219000736428262 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_102 (.en(wire_76), .in(wire_140), .out(wire_54_8));
  TC_LessU # (.UUID(64'd70784060852193480 ^ UUID), .BIT_WIDTH(64'd16)) LessU16_103 (.in0(wire_35), .in1(wire_97), .out(wire_140));
  TC_Or # (.UUID(64'd2633850717105506955 ^ UUID), .BIT_WIDTH(64'd1)) Or_104 (.in0(wire_140), .in1(wire_197), .out(wire_70));
  TC_Not # (.UUID(64'd2994142474806724920 ^ UUID), .BIT_WIDTH(64'd1)) Not_105 (.in(wire_197), .out(wire_206));
  TC_Equal # (.UUID(64'd4180772301230732474 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_106 (.in0(wire_97), .in1(wire_35), .out(wire_197));
  TC_LessU # (.UUID(64'd3216607671565821129 ^ UUID), .BIT_WIDTH(64'd16)) LessU16_107 (.in0(wire_97), .in1(wire_35), .out(wire_107));
  TC_Or # (.UUID(64'd1733367887190953979 ^ UUID), .BIT_WIDTH(64'd1)) Or_108 (.in0(wire_197), .in1(wire_107), .out(wire_243));
  TC_Equal # (.UUID(64'd2756161344151621510 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_109 (.in0({{8{1'b0}}, wire_398 }), .in1(wire_97), .out(wire_93));
  TC_Constant # (.UUID(64'd14059539423913175 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h0)) Constant8_110 (.out(wire_398));
  TC_Not # (.UUID(64'd2912282656104074477 ^ UUID), .BIT_WIDTH(64'd1)) Not_111 (.in(wire_93), .out(wire_299));
  TC_Switch # (.UUID(64'd338503895939097385 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_112 (.en(wire_192), .in(wire_93), .out(wire_54_2));
  TC_Switch # (.UUID(64'd2974250978505416008 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_113 (.en(wire_40), .in(wire_97), .out(wire_28));
  TC_Switch # (.UUID(64'd294942412853573551 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_114 (.en(wire_11), .in(wire_46), .out(wire_127_0));
  TC_Switch # (.UUID(64'd2530020128287448865 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_115 (.en(wire_260), .in(wire_84), .out(wire_127_1));
  TC_Not # (.UUID(64'd1944022449022311076 ^ UUID), .BIT_WIDTH(64'd1)) Not_116 (.in(wire_11), .out(wire_260));
  TC_Switch # (.UUID(64'd640117511591385720 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_117 (.en(wire_338), .in(wire_97), .out(wire_1_7[15:0]));
  TC_Clock # (.UUID(64'd473244454118914110 ^ UUID)) Clock_118 (.clk(clk), .rst(rst), .out(wire_11));
  TC_Switch # (.UUID(64'd3240978896697767469 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_119 (.en(wire_105), .in(wire_105), .out(wire_54_5));
  TC_Mux # (.UUID(64'd4327728578462997473 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_120 (.sel(wire_47), .in0(wire_74), .in1(wire_283), .out(wire_84));
  TC_Not # (.UUID(64'd2335834251709147674 ^ UUID), .BIT_WIDTH(64'd1)) Not_121 (.in(wire_212), .out(wire_298));
  TC_Switch # (.UUID(64'd1177966569030928993 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_122 (.en(wire_212), .in(wire_136), .out(wire_1_4[15:0]));
  TC_Switch # (.UUID(64'd4085565154656183842 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_123 (.en(wire_95), .in(wire_403), .out(wire_1_0[15:0]));
  TC_IndexerByte # (.UUID(64'd82359665637793120 ^ UUID), .INDEX(64'd2)) IndexerByte_124 (.in({{32{1'b0}}, wire_139 }), .out(wire_373));
  TC_Switch # (.UUID(64'd691486037870060392 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_125 (.en(wire_226), .in(wire_132), .out(wire_43));
  TC_IndexerBit # (.UUID(64'd1630189301439907508 ^ UUID), .INDEX(64'd4)) IndexerBit_126 (.in({{56{1'b0}}, wire_34 }), .out(wire_5));
  TC_IndexerBit # (.UUID(64'd2208263359456905046 ^ UUID), .INDEX(64'd5)) IndexerBit_127 (.in({{56{1'b0}}, wire_34 }), .out(wire_55));
  TC_IndexerByte # (.UUID(64'd2160584388702904456 ^ UUID), .INDEX(64'd3)) IndexerByte_128 (.in({{32{1'b0}}, wire_139 }), .out(wire_34));
  TC_Not # (.UUID(64'd904891828379418593 ^ UUID), .BIT_WIDTH(64'd1)) Not_129 (.in(wire_55), .out(wire_301));
  TC_Constant # (.UUID(64'd3538634162844758805 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hFF)) Constant8_130 (.out(wire_293));
  TC_Constant # (.UUID(64'd2648359173322761393 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hFE)) Constant8_131 (.out(wire_116));
  TC_Maker16 # (.UUID(64'd4168581648613032575 ^ UUID)) Maker16_132 (.in0(wire_293), .in1(wire_116), .out(wire_407));
  TC_Mux # (.UUID(64'd3090540701337537666 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_133 (.sel(wire_49), .in0(wire_239), .in1(wire_283), .out(wire_46));
  TC_Maker16 # (.UUID(64'd851087207377417069 ^ UUID)) Maker16_134 (.in0(wire_274), .in1(wire_6), .out(wire_307));
  TC_Constant # (.UUID(64'd381873739773538407 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hFF)) Constant8_135 (.out(wire_274));
  TC_Mux # (.UUID(64'd4592224200207251913 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_136 (.sel(wire_301), .in0(wire_172), .in1(wire_263), .out(wire_149));
  TC_Equal # (.UUID(64'd3099658865939077738 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_137 (.in0(wire_43), .in1(16'd0), .out(wire_267));
  TC_Not # (.UUID(64'd4471125710935676612 ^ UUID), .BIT_WIDTH(64'd1)) Not_138 (.in(wire_267), .out(wire_186));
  TC_IndexerBit # (.UUID(64'd460606693629125729 ^ UUID), .INDEX(64'd4)) IndexerBit_139 (.in({{56{1'b0}}, wire_110 }), .out(wire_207));
  TC_IndexerBit # (.UUID(64'd1499309531990315318 ^ UUID), .INDEX(64'd1)) IndexerBit_140 (.in({{56{1'b0}}, wire_110 }), .out(wire_227));
  TC_Or3 # (.UUID(64'd3834216222200410896 ^ UUID), .BIT_WIDTH(64'd1)) Or3_141 (.in0(wire_75), .in1(wire_358), .in2(wire_319), .out(wire_40));
  TC_IndexerBit # (.UUID(64'd345801079655292532 ^ UUID), .INDEX(64'd2)) IndexerBit_142 (.in({{56{1'b0}}, wire_110 }), .out(wire_358));
  TC_IndexerBit # (.UUID(64'd3857678701898454921 ^ UUID), .INDEX(64'd3)) IndexerBit_143 (.in({{56{1'b0}}, wire_110 }), .out(wire_75));
  TC_IndexerBit # (.UUID(64'd1094550749412879412 ^ UUID), .INDEX(64'd5)) IndexerBit_144 (.in({{56{1'b0}}, wire_110 }), .out(wire_0));
  TC_Not # (.UUID(64'd295801019876953925 ^ UUID), .BIT_WIDTH(64'd1)) Not_145 (.in(wire_334), .out(wire_120));
  TC_Equal # (.UUID(64'd3140328761418953014 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_146 (.in0(wire_46), .in1(16'd0), .out(wire_396));
  TC_Not # (.UUID(64'd4400946405007906585 ^ UUID), .BIT_WIDTH(64'd1)) Not_147 (.in(wire_394), .out(wire_156));
  TC_IndexerByte # (.UUID(64'd2633087214037843825 ^ UUID), .INDEX(64'd3)) IndexerByte_148 (.in({{32{1'b0}}, wire_139 }), .out(wire_110));
  TC_Equal # (.UUID(64'd2561182539117830921 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_149 (.in0(16'd0), .in1(wire_84), .out(wire_394));
  TC_IndexerBit # (.UUID(64'd2047893359182210890 ^ UUID), .INDEX(64'd0)) IndexerBit_150 (.in(wire_10), .out(wire_14));
  TC_IndexerBit # (.UUID(64'd3859884203355858265 ^ UUID), .INDEX(64'd1)) IndexerBit_151 (.in(wire_10), .out(wire_99));
  TC_IndexerBit # (.UUID(64'd4287739567158645737 ^ UUID), .INDEX(64'd2)) IndexerBit_152 (.in(wire_10), .out(wire_25));
  TC_IndexerBit # (.UUID(64'd777253982648504148 ^ UUID), .INDEX(64'd3)) IndexerBit_153 (.in(wire_10), .out(wire_21));
  TC_IndexerBit # (.UUID(64'd1771789865896455183 ^ UUID), .INDEX(64'd4)) IndexerBit_154 (.in(wire_10), .out(wire_213));
  TC_IndexerBit # (.UUID(64'd3105812192345802732 ^ UUID), .INDEX(64'd6)) IndexerBit_155 (.in(wire_10), .out(wire_18));
  TC_IndexerBit # (.UUID(64'd3077471030622112266 ^ UUID), .INDEX(64'd7)) IndexerBit_156 (.in(wire_10), .out(wire_114));
  TC_Not # (.UUID(64'd2159748274689718655 ^ UUID), .BIT_WIDTH(64'd1)) Not_157 (.in(wire_396), .out(wire_367));
  TC_Splitter16 # (.UUID(64'd1069070463351244943 ^ UUID)) Splitter16_158 (.in(wire_10[15:0]), .out0(), .out1(wire_150));
  TC_Switch # (.UUID(64'd3542778498052595836 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_159 (.en(wire_146), .in(wire_381[15:0]), .out(wire_1_20[15:0]));
  TC_Not # (.UUID(64'd944680686405816927 ^ UUID), .BIT_WIDTH(64'd1)) Not_160 (.in(wire_183), .out(wire_316));
  TC_Switch # (.UUID(64'd816465745217087424 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_161 (.en(wire_229), .in(wire_35), .out(wire_15));
  TC_Switch # (.UUID(64'd209623535459112064 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_162 (.en(wire_229), .in(wire_97), .out(wire_189));
  TC_And # (.UUID(64'd2522855677877010919 ^ UUID), .BIT_WIDTH(64'd1)) And_163 (.in0(wire_229), .in1(wire_12), .out(wire_146));
  TC_Equal # (.UUID(64'd2756262866884777429 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_164 (.in0(8'd0), .in1(wire_189[7:0]), .out(wire_12));
  TC_Equal # (.UUID(64'd1714264829042601315 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_165 (.in0(wire_150), .in1(wire_134), .out(wire_229));
  TC_Constant # (.UUID(64'd2907468583675662890 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_166 (.out(wire_134));
  TC_Mux # (.UUID(64'd2441497898305995710 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_167 (.sel(wire_5), .in0(wire_161), .in1(wire_172), .out(wire_239));
  TC_Switch # (.UUID(64'd3809517357945142409 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_168 (.en(wire_214), .in(wire_126[15:0]), .out(wire_167));
  TC_Not # (.UUID(64'd4003951151984714090 ^ UUID), .BIT_WIDTH(64'd1)) Not_169 (.in(wire_114), .out(wire_311));
  TC_IndexerBit # (.UUID(64'd1553590145675495351 ^ UUID), .INDEX(64'd5)) IndexerBit_170 (.in(wire_10), .out(wire_212));
  TC_Not # (.UUID(64'd3312304652180753239 ^ UUID), .BIT_WIDTH(64'd1)) Not_171 (.in(wire_18), .out(wire_226));
  TC_Constant # (.UUID(64'd2729531845625831067 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_172 (.out(wire_236));
  TC_Not # (.UUID(64'd2538698523318428916 ^ UUID), .BIT_WIDTH(64'd1)) Not_173 (.in(wire_339), .out(wire_329));
  TC_Constant # (.UUID(64'd2179489257373318160 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_174 (.out(wire_122));
  TC_Mux # (.UUID(64'd2429066787419951843 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_175 (.sel(wire_4), .in0(wire_35), .in1({{8{1'b0}}, wire_122 }), .out(wire_62));
  TC_Switch # (.UUID(64'd391371808230282023 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_176 (.en(wire_209), .in(wire_345), .out(wire_357));
  TC_Constant # (.UUID(64'd2691125905525222303 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1F)) Constant8_177 (.out(wire_390));
  TC_IndexerByte # (.UUID(64'd2112170900386343144 ^ UUID), .INDEX(64'd3)) IndexerByte_178 (.in({{32{1'b0}}, wire_139 }), .out(wire_328));
  TC_IndexerBit # (.UUID(64'd2727080739164391000 ^ UUID), .INDEX(64'd6)) IndexerBit_179 (.in({{56{1'b0}}, wire_328 }), .out(wire_255));
  TC_Switch # (.UUID(64'd2160087561000370162 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_180 (.en(wire_255), .in(wire_255), .out(wire_54_9));
  TC_Switch # (.UUID(64'd592302940647155691 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_181 (.en(wire_222), .in({{15{1'b0}}, wire_364 }), .out(wire_1_11[15:0]));
  TC_Or # (.UUID(64'd3278179513885088927 ^ UUID), .BIT_WIDTH(64'd1)) Or_182 (.in0(wire_222), .in1(wire_113), .out(wire_230));
  TC_Equal # (.UUID(64'd4033274235037801114 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_183 (.in0(wire_346), .in1(wire_348), .out(wire_222));
  TC_Not # (.UUID(64'd1697593568395826930 ^ UUID), .BIT_WIDTH(64'd1)) Not_184 (.in(wire_113), .out(wire_372));
  TC_Splitter16 # (.UUID(64'd962308306064647197 ^ UUID)) Splitter16_185 (.in(wire_10[15:0]), .out0(), .out1(wire_346));
  TC_Constant # (.UUID(64'd3037869375563223000 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h2)) Constant8_186 (.out(wire_348));
  TC_DelayLine # (.UUID(64'd4275385609773382257 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_187 (.clk(clk), .rst(rst), .in(wire_32), .out(wire_113));
  TC_Switch # (.UUID(64'd1286392688347840013 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_188 (.en(wire_372), .in(wire_230), .out(wire_32));
  TC_Splitter16 # (.UUID(64'd815166994044352782 ^ UUID)) Splitter16_189 (.in(wire_10[15:0]), .out0(), .out1(wire_340));
  TC_IndexerByte # (.UUID(64'd4056757385308142069 ^ UUID), .INDEX(64'd1)) IndexerByte_190 (.in(wire_169), .out(wire_275));
  TC_IndexerByte # (.UUID(64'd4445007758314830950 ^ UUID), .INDEX(64'd0)) IndexerByte_191 (.in(wire_169), .out(wire_168));
  TC_Maker16 # (.UUID(64'd1879612468053834457 ^ UUID)) Maker16_192 (.in0(wire_168), .in1(wire_275), .out(wire_152));
  TC_Switch # (.UUID(64'd220823607166135876 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_193 (.en(wire_237), .in(wire_152), .out(wire_1_15[15:0]));
  TC_Equal # (.UUID(64'd3724760983101447498 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_194 (.in0(wire_340), .in1(wire_291), .out(wire_237));
  TC_Constant # (.UUID(64'd1337227511337026411 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h3)) Constant8_195 (.out(wire_291));
  TC_Timing # (.UUID(64'd2799049267103079424 ^ UUID)) Timing_196 (.en(wire_237), .out(wire_169));
  TC_Program # (.UUID(64'd3721980137216604240 ^ UUID), .WORD_WIDTH(64'd8), .DEFAULT_FILE_NAME("Program_33A7213703DAF850.w8.bin"), .ARG_SIG("Program_33A7213703DAF850=%s")) Program_197 (.clk(clk), .rst(rst), .address(wire_97), .out0(wire_187), .out1(), .out2(), .out3());
  TC_Splitter16 # (.UUID(64'd4461787469973933422 ^ UUID)) Splitter16_198 (.in(wire_10[15:0]), .out0(), .out1(wire_123));
  TC_Equal # (.UUID(64'd1988770091565985332 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_199 (.in0(wire_123), .in1(wire_106), .out(wire_268));
  TC_Constant # (.UUID(64'd2565543928344869306 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h5)) Constant8_200 (.out(wire_106));
  TC_Switch # (.UUID(64'd4105771623231641306 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_201 (.en(wire_268), .in(wire_187[15:0]), .out(wire_1_18[15:0]));
  TC_Equal # (.UUID(64'd551722571517782638 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_202 (.in0(16'd0), .in1(wire_189), .out(wire_183));
  TC_Register # (.UUID(64'd4364107987795409853 ^ UUID), .BIT_WIDTH(64'd16)) Register16_203 (.clk(clk), .rst(rst), .load(wire_277), .save(wire_277), .in(wire_235), .out(wire_85));
  TC_Constant # (.UUID(64'd1415884859697557611 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_204 (.out(wire_173));
  TC_IndexerBit # (.UUID(64'd535377880148297947 ^ UUID), .INDEX(64'd3)) IndexerBit_205 (.in({{56{1'b0}}, wire_34 }), .out(wire_47));
  TC_Register # (.UUID(64'd2160598746671012754 ^ UUID), .BIT_WIDTH(64'd16)) Register16_206 (.clk(clk), .rst(rst), .load(wire_105), .save(wire_105), .in(wire_45), .out(wire_8));
  TC_Add # (.UUID(64'd1442806402229030427 ^ UUID), .BIT_WIDTH(64'd16)) Add16_207 (.in0(wire_400), .in1(wire_407), .ci(1'd0), .out(wire_172), .co());
  TC_Or # (.UUID(64'd2188959817660993009 ^ UUID), .BIT_WIDTH(64'd1)) Or_208 (.in0(wire_5), .in1(wire_55), .out(wire_105));
  TC_IndexerBit # (.UUID(64'd3588176080026118662 ^ UUID), .INDEX(64'd2)) IndexerBit_209 (.in({{56{1'b0}}, wire_34 }), .out(wire_49));
  TC_Mux # (.UUID(64'd4063471477342436371 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_210 (.sel(wire_55), .in0(wire_388), .in1(wire_8), .out(wire_400));
  TC_Mux # (.UUID(64'd527759690959107192 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_211 (.sel(wire_47), .in0(wire_285), .in1(wire_85), .out(wire_185));
  TC_Switch # (.UUID(64'd1362725833065582892 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_212 (.en(wire_49), .in(wire_235), .out(wire_285));
  TC_Switch # (.UUID(64'd1756831740426205013 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_213 (.en(wire_5), .in(wire_45), .out(wire_388));
  TC_Add # (.UUID(64'd2930665708224337659 ^ UUID), .BIT_WIDTH(64'd16)) Add16_214 (.in0(wire_85), .in1(wire_204), .ci(1'd0), .out(wire_235), .co());
  TC_Constant # (.UUID(64'd3137150186803814383 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hF0)) Constant8_215 (.out(wire_6));
  TC_Add # (.UUID(64'd432537638553101254 ^ UUID), .BIT_WIDTH(64'd16)) Add16_216 (.in0(wire_8), .in1(wire_336), .ci(1'd0), .out(wire_45), .co());
  TC_IndexerBit # (.UUID(64'd561707948535025464 ^ UUID), .INDEX(64'd4)) IndexerBit_217 (.in({{56{1'b0}}, wire_34 }), .out(wire_397));
  TC_Constant # (.UUID(64'd1695694096694981758 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_218 (.out(wire_89));
  TC_IndexerBit # (.UUID(64'd2331812482237933900 ^ UUID), .INDEX(64'd0)) IndexerBit_219 (.in({{56{1'b0}}, wire_96 }), .out(wire_319));
  TC_Neg # (.UUID(64'd1821476619534246961 ^ UUID), .BIT_WIDTH(64'd16)) Neg16_220 (.in({{8{1'b0}}, wire_89 }), .out(wire_401));
  TC_Mux # (.UUID(64'd1539425850473868597 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_221 (.sel(wire_397), .in0(wire_401), .in1({{8{1'b0}}, wire_89 }), .out(wire_336));
  TC_Mux # (.UUID(64'd3572805427243657698 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_222 (.sel(wire_49), .in0(wire_286), .in1({{8{1'b0}}, wire_173 }), .out(wire_204));
  TC_Neg # (.UUID(64'd2090057048615449572 ^ UUID), .BIT_WIDTH(64'd16)) Neg16_223 (.in({{8{1'b0}}, wire_173 }), .out(wire_286));
  TC_IOSwitch # (.UUID(64'd2846053541171193881 ^ UUID), .BIT_WIDTH(64'd8)) LevelOutputArch_224 (.in(wire_97[7:0]), .en(wire_92), .out(arch_output_value));
  TC_Switch # (.UUID(64'd210661621448949326 ^ UUID), .BIT_WIDTH(64'd8)) LevelInputArch_225 (.en(wire_335), .in(arch_input_value), .out(wire_1_19[7:0]));
  TC_Splitter16 # (.UUID(64'd2775342692045340835 ^ UUID)) Splitter16_226 (.in(wire_10[15:0]), .out0(), .out1(wire_57));
  TC_Equal # (.UUID(64'd4532639728004948159 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_227 (.in0(wire_57), .in1(wire_208), .out(wire_224));
  TC_Equal # (.UUID(64'd3745587913460272427 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_228 (.in0(wire_399), .in1(wire_57), .out(wire_59));
  TC_Constant # (.UUID(64'd951998662890801082 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6)) Constant8_229 (.out(wire_399));
  TC_Constant # (.UUID(64'd2262634952183580731 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7)) Constant8_230 (.out(wire_208));
  TC_Switch # (.UUID(64'd1419008802292368204 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_231 (.en(wire_300), .in(wire_59), .out(wire_335));
  TC_Clock # (.UUID(64'd150335021447124340 ^ UUID)) Clock_232 (.clk(clk), .rst(rst), .out(wire_300));
  TC_Switch # (.UUID(64'd3781955660154943019 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_233 (.en(wire_391), .in(wire_224), .out(wire_92));
  TC_Not # (.UUID(64'd248590985388437467 ^ UUID), .BIT_WIDTH(64'd1)) Not_234 (.in(wire_300), .out(wire_391));
  TC_RamDualLoad # (.UUID(64'd1162091816344660036 ^ UUID), .WORD_WIDTH(64'd16), .WORD_COUNT(64'd65536)) RamDualLoad_235 (.clk(clk), .rst(rst), .load0(wire_156), .save(wire_367), .address0({{16{1'b0}}, wire_127 }), .in({{48{1'b0}}, wire_179 }), .load1(wire_186), .address1({{16{1'b0}}, wire_43 }), .out0(wire_379), .out1(wire_218));
  TC_Ram # (.UUID(64'd2071862132571227302 ^ UUID), .WORD_WIDTH(64'd16), .WORD_COUNT(64'd65536)) Ram_236 (.clk(clk), .rst(rst), .load(wire_183), .save(wire_316), .address({{16{1'b0}}, wire_15 }), .in0({{48{1'b0}}, wire_189 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_381), .out1(), .out2(), .out3());
  TC_FileLoader # (.UUID(64'd1149854990232492044 ^ UUID), .DEFAULT_FILE_NAME("image.dat")) FileLoader_237 (.clk(clk), .rst(rst), .en(wire_182), .address({{48{1'b0}}, wire_97 }), .out(wire_1_13));
  TC_Splitter16 # (.UUID(64'd2684349980131024015 ^ UUID)) Splitter16_238 (.in(wire_10[15:0]), .out0(), .out1(wire_141));
  TC_Equal # (.UUID(64'd4369488988257915881 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_239 (.in0(wire_141), .in1(wire_137), .out(wire_182));
  TC_Constant # (.UUID(64'd3823619217162964047 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h8)) Constant8_240 (.out(wire_137));
  TC_Ror # (.UUID(64'd445352019034615982 ^ UUID), .BIT_WIDTH(64'd16)) Ror16_241 (.in(wire_97), .shift(wire_35[7:0]), .out(wire_147));
  TC_DotMatrixDisplay # (.UUID(64'd4586922663638092405 ^ UUID)) DotMatrixDisplay_242 (.clk(clk), .rst(rst), .en_y(wire_219[0:0]), .en_x(wire_165[0:0]), .color_info(wire_219), .pixel_info(wire_165));
  TC_DotMatrixDisplay # (.UUID(64'd768543756621643271 ^ UUID)) DotMatrixDisplay_243 (.clk(clk), .rst(rst), .en_y(wire_101[0:0]), .en_x(wire_165[0:0]), .color_info(wire_101), .pixel_info(wire_165));
  TC_DotMatrixDisplay # (.UUID(64'd1312987478703542956 ^ UUID)) DotMatrixDisplay_244 (.clk(clk), .rst(rst), .en_y(wire_244[0:0]), .en_x(wire_165[0:0]), .color_info(wire_244), .pixel_info(wire_165));
  TC_DotMatrixDisplay # (.UUID(64'd3831511369089243381 ^ UUID)) DotMatrixDisplay_245 (.clk(clk), .rst(rst), .en_y(wire_56[0:0]), .en_x(wire_165[0:0]), .color_info(wire_56), .pixel_info(wire_165));
  TC_DotMatrixDisplay # (.UUID(64'd544763639986031707 ^ UUID)) DotMatrixDisplay_246 (.clk(clk), .rst(rst), .en_y(wire_178[0:0]), .en_x(wire_165[0:0]), .color_info(wire_178), .pixel_info(wire_165));
  TC_DotMatrixDisplay # (.UUID(64'd2831844111636891909 ^ UUID)) DotMatrixDisplay_247 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_165[0:0]), .color_info(wire_22), .pixel_info(wire_165));
  TC_DotMatrixDisplay # (.UUID(64'd803399427566320925 ^ UUID)) DotMatrixDisplay_248 (.clk(clk), .rst(rst), .en_y(wire_219[0:0]), .en_x(wire_191[0:0]), .color_info(wire_219), .pixel_info(wire_191));
  TC_DotMatrixDisplay # (.UUID(64'd3855072706384208530 ^ UUID)) DotMatrixDisplay_249 (.clk(clk), .rst(rst), .en_y(wire_101[0:0]), .en_x(wire_191[0:0]), .color_info(wire_101), .pixel_info(wire_191));
  TC_DotMatrixDisplay # (.UUID(64'd4206739403808363797 ^ UUID)) DotMatrixDisplay_250 (.clk(clk), .rst(rst), .en_y(wire_244[0:0]), .en_x(wire_191[0:0]), .color_info(wire_244), .pixel_info(wire_191));
  TC_DotMatrixDisplay # (.UUID(64'd1651693078729037187 ^ UUID)) DotMatrixDisplay_251 (.clk(clk), .rst(rst), .en_y(wire_56[0:0]), .en_x(wire_191[0:0]), .color_info(wire_56), .pixel_info(wire_191));
  TC_DotMatrixDisplay # (.UUID(64'd866725564843264959 ^ UUID)) DotMatrixDisplay_252 (.clk(clk), .rst(rst), .en_y(wire_178[0:0]), .en_x(wire_191[0:0]), .color_info(wire_178), .pixel_info(wire_191));
  TC_DotMatrixDisplay # (.UUID(64'd1713126292273528914 ^ UUID)) DotMatrixDisplay_253 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_191[0:0]), .color_info(wire_22), .pixel_info(wire_191));
  TC_DotMatrixDisplay # (.UUID(64'd464335165834344681 ^ UUID)) DotMatrixDisplay_254 (.clk(clk), .rst(rst), .en_y(wire_219[0:0]), .en_x(wire_19[0:0]), .color_info(wire_219), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd212104235248741642 ^ UUID)) DotMatrixDisplay_255 (.clk(clk), .rst(rst), .en_y(wire_101[0:0]), .en_x(wire_19[0:0]), .color_info(wire_101), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd4116412079736924536 ^ UUID)) DotMatrixDisplay_256 (.clk(clk), .rst(rst), .en_y(wire_244[0:0]), .en_x(wire_19[0:0]), .color_info(wire_244), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd3195163277462157351 ^ UUID)) DotMatrixDisplay_257 (.clk(clk), .rst(rst), .en_y(wire_56[0:0]), .en_x(wire_19[0:0]), .color_info(wire_56), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd2373424346728527832 ^ UUID)) DotMatrixDisplay_258 (.clk(clk), .rst(rst), .en_y(wire_178[0:0]), .en_x(wire_19[0:0]), .color_info(wire_178), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd4464466339432778604 ^ UUID)) DotMatrixDisplay_259 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_19[0:0]), .color_info(wire_22), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd1989401320784160937 ^ UUID)) DotMatrixDisplay_260 (.clk(clk), .rst(rst), .en_y(wire_219[0:0]), .en_x(wire_50[0:0]), .color_info(wire_219), .pixel_info(wire_50));
  TC_DotMatrixDisplay # (.UUID(64'd4346815494554460150 ^ UUID)) DotMatrixDisplay_261 (.clk(clk), .rst(rst), .en_y(wire_56[0:0]), .en_x(wire_50[0:0]), .color_info(wire_56), .pixel_info(wire_50));
  TC_DotMatrixDisplay # (.UUID(64'd4448216468649510302 ^ UUID)) DotMatrixDisplay_262 (.clk(clk), .rst(rst), .en_y(wire_178[0:0]), .en_x(wire_50[0:0]), .color_info(wire_178), .pixel_info(wire_50));
  TC_DotMatrixDisplay # (.UUID(64'd2608578660833632206 ^ UUID)) DotMatrixDisplay_263 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_50[0:0]), .color_info(wire_22), .pixel_info(wire_50));
  TC_Or # (.UUID(64'd2774518916655491254 ^ UUID), .BIT_WIDTH(64'd32)) Or32_264 (.in0({{31{1'b0}}, wire_170 }), .in1(wire_9), .out(wire_219));
  TC_Or # (.UUID(64'd3577024797358561642 ^ UUID), .BIT_WIDTH(64'd32)) Or32_265 (.in0({{31{1'b0}}, wire_65 }), .in1(wire_9), .out(wire_101));
  TC_Or # (.UUID(64'd2364218693127516361 ^ UUID), .BIT_WIDTH(64'd32)) Or32_266 (.in0({{31{1'b0}}, wire_216 }), .in1(wire_9), .out(wire_56));
  TC_Or # (.UUID(64'd4211847430470965668 ^ UUID), .BIT_WIDTH(64'd32)) Or32_267 (.in0({{31{1'b0}}, wire_355 }), .in1(wire_9), .out(wire_178));
  TC_Or # (.UUID(64'd3856510800564153436 ^ UUID), .BIT_WIDTH(64'd32)) Or32_268 (.in0({{31{1'b0}}, wire_121 }), .in1(wire_9), .out(wire_22));
  TC_Decoder3 # (.UUID(64'd345945806527240068 ^ UUID)) Decoder3_269 (.dis(1'd0), .sel0(wire_7), .sel1(wire_408), .sel2(wire_118), .out0(wire_170), .out1(wire_65), .out2(wire_276), .out3(wire_216), .out4(wire_355), .out5(wire_121), .out6(), .out7());
  TC_Or # (.UUID(64'd1220236455381113553 ^ UUID), .BIT_WIDTH(64'd64)) Or64_270 (.in0(wire_63), .in1({{63{1'b0}}, wire_343 }), .out(wire_250));
  TC_Or # (.UUID(64'd4088311446664524645 ^ UUID), .BIT_WIDTH(64'd64)) Or64_271 (.in0(wire_63), .in1({{63{1'b0}}, wire_166 }), .out(wire_290));
  TC_Or # (.UUID(64'd4495256993990392420 ^ UUID), .BIT_WIDTH(64'd64)) Or64_272 (.in0(wire_63), .in1({{63{1'b0}}, wire_61 }), .out(wire_386));
  TC_Decoder2 # (.UUID(64'd1792850179932055927 ^ UUID)) Decoder2_273 (.sel0(wire_258), .sel1(wire_164), .out0(wire_343), .out1(wire_166), .out2(wire_314), .out3(wire_61));
  TC_Or # (.UUID(64'd2399075346851224651 ^ UUID), .BIT_WIDTH(64'd64)) Or64_274 (.in0(wire_63), .in1({{63{1'b0}}, wire_314 }), .out(wire_248));
  TC_Or # (.UUID(64'd1701960925663082587 ^ UUID), .BIT_WIDTH(64'd64)) Or64_275 (.in0(wire_248), .in1(wire_217), .out(wire_19));
  TC_Or # (.UUID(64'd2764878805242022165 ^ UUID), .BIT_WIDTH(64'd64)) Or64_276 (.in0(wire_386), .in1(wire_217), .out(wire_50));
  TC_Or # (.UUID(64'd2748551646898479399 ^ UUID), .BIT_WIDTH(64'd64)) Or64_277 (.in0(wire_290), .in1(wire_217), .out(wire_191));
  TC_Or # (.UUID(64'd579758728963367249 ^ UUID), .BIT_WIDTH(64'd64)) Or64_278 (.in0(wire_250), .in1(wire_217), .out(wire_165));
  TC_IndexerBit # (.UUID(64'd1915715909516237622 ^ UUID), .INDEX(64'd0)) IndexerBit_279 (.in({{48{1'b0}}, wire_39 }), .out(wire_7));
  TC_IndexerBit # (.UUID(64'd384185582563507733 ^ UUID), .INDEX(64'd1)) IndexerBit_280 (.in({{48{1'b0}}, wire_39 }), .out(wire_408));
  TC_IndexerBit # (.UUID(64'd1844140052021087840 ^ UUID), .INDEX(64'd2)) IndexerBit_281 (.in({{48{1'b0}}, wire_39 }), .out(wire_118));
  TC_Or # (.UUID(64'd2562615352787499523 ^ UUID), .BIT_WIDTH(64'd32)) Or32_282 (.in0({{31{1'b0}}, wire_276 }), .in1(wire_9), .out(wire_244));
  TC_DotMatrixDisplay # (.UUID(64'd1877295406034505077 ^ UUID)) DotMatrixDisplay_283 (.clk(clk), .rst(rst), .en_y(wire_244[0:0]), .en_x(wire_50[0:0]), .color_info(wire_244), .pixel_info(wire_50));
  TC_DotMatrixDisplay # (.UUID(64'd3592707041588415280 ^ UUID)) DotMatrixDisplay_284 (.clk(clk), .rst(rst), .en_y(wire_101[0:0]), .en_x(wire_50[0:0]), .color_info(wire_101), .pixel_info(wire_50));
  TC_IndexerBit # (.UUID(64'd1397832739463884705 ^ UUID), .INDEX(64'd1)) IndexerBit_285 (.in({{56{1'b0}}, wire_228 }), .out(wire_164));
  TC_Constant # (.UUID(64'd370664463030471557 ^ UUID), .BIT_WIDTH(64'd64), .value(64'h100000000000000)) Constant64_286 (.out(wire_217));
  TC_Maker8 # (.UUID(64'd2588821264127475169 ^ UUID)) Maker8_287 (.in0(wire_103), .in1(wire_72), .in2(wire_103), .in3(wire_72), .in4(wire_103), .in5(wire_72), .in6(wire_103), .in7(wire_72), .out(wire_100));
  TC_Maker8 # (.UUID(64'd2828170759771675122 ^ UUID)) Maker8_288 (.in0(wire_37), .in1(wire_33), .in2(wire_37), .in3(wire_33), .in4(wire_37), .in5(wire_33), .in6(wire_37), .in7(wire_33), .out(wire_225));
  TC_Maker8 # (.UUID(64'd2415308843918290587 ^ UUID)) Maker8_289 (.in0(wire_24), .in1(wire_259), .in2(wire_24), .in3(wire_259), .in4(wire_24), .in5(wire_259), .in6(wire_24), .in7(wire_259), .out(wire_241));
  TC_IndexerBit # (.UUID(64'd1843601702595912724 ^ UUID), .INDEX(64'd6)) IndexerBit_290 (.in({{56{1'b0}}, wire_68 }), .out(wire_103));
  TC_IndexerBit # (.UUID(64'd3753608481866364619 ^ UUID), .INDEX(64'd7)) IndexerBit_291 (.in({{56{1'b0}}, wire_68 }), .out(wire_72));
  TC_IndexerBit # (.UUID(64'd4255822523224537977 ^ UUID), .INDEX(64'd4)) IndexerBit_292 (.in({{56{1'b0}}, wire_68 }), .out(wire_37));
  TC_IndexerBit # (.UUID(64'd933032544826559249 ^ UUID), .INDEX(64'd5)) IndexerBit_293 (.in({{56{1'b0}}, wire_68 }), .out(wire_33));
  TC_IndexerBit # (.UUID(64'd4120795911758374986 ^ UUID), .INDEX(64'd2)) IndexerBit_294 (.in({{56{1'b0}}, wire_68 }), .out(wire_24));
  TC_IndexerBit # (.UUID(64'd3957574907750575317 ^ UUID), .INDEX(64'd3)) IndexerBit_295 (.in({{56{1'b0}}, wire_68 }), .out(wire_259));
  TC_IndexerBit # (.UUID(64'd630305000696767227 ^ UUID), .INDEX(64'd0)) IndexerBit_296 (.in({{56{1'b0}}, wire_228 }), .out(wire_258));
  TC_IndexerByte # (.UUID(64'd2466525370095194356 ^ UUID), .INDEX(64'd1)) IndexerByte_297 (.in({{48{1'b0}}, wire_39 }), .out(wire_228));
  TC_Maker32 # (.UUID(64'd3137312401582712707 ^ UUID)) Maker32_298 (.in0(8'd0), .in1(wire_241), .in2(wire_225), .in3(wire_100), .out(wire_9));
  TC_Maker8 # (.UUID(64'd849915623509302596 ^ UUID)) Maker8_299 (.in0(wire_196), .in1(wire_234), .in2(wire_2), .in3(wire_289), .in4(wire_90), .in5(wire_252), .in6(wire_223), .in7(wire_245), .out(wire_131));
  TC_Maker8 # (.UUID(64'd1347595989490070695 ^ UUID)) Maker8_300 (.in0(wire_409), .in1(wire_254), .in2(wire_406), .in3(wire_371), .in4(wire_112), .in5(wire_310), .in6(wire_342), .in7(wire_73), .out(wire_304));
  TC_Decoder3 # (.UUID(64'd2440547940564590289 ^ UUID)) Decoder3_301 (.dis(wire_279), .sel0(wire_23), .sel1(wire_138), .sel2(wire_30), .out0(wire_196), .out1(wire_234), .out2(wire_2), .out3(wire_289), .out4(wire_90), .out5(wire_252), .out6(wire_223), .out7(wire_245));
  TC_Decoder3 # (.UUID(64'd2079858873611333618 ^ UUID)) Decoder3_302 (.dis(wire_374), .sel0(wire_23), .sel1(wire_138), .sel2(wire_30), .out0(wire_409), .out1(wire_254), .out2(wire_406), .out3(wire_371), .out4(wire_112), .out5(wire_310), .out6(wire_342), .out7(wire_73));
  TC_Maker8 # (.UUID(64'd3108610901977927566 ^ UUID)) Maker8_303 (.in0(wire_321), .in1(wire_69), .in2(wire_330), .in3(wire_36), .in4(wire_180), .in5(wire_48), .in6(wire_395), .in7(wire_272), .out(wire_256));
  TC_Decoder3 # (.UUID(64'd1913239957499811182 ^ UUID)) Decoder3_304 (.dis(wire_201), .sel0(wire_23), .sel1(wire_138), .sel2(wire_30), .out0(wire_321), .out1(wire_69), .out2(wire_330), .out3(wire_36), .out4(wire_180), .out5(wire_48), .out6(wire_395), .out7(wire_272));
  TC_IndexerBit # (.UUID(64'd2823428697791387290 ^ UUID), .INDEX(64'd3)) IndexerBit_305 (.in({{56{1'b0}}, wire_71 }), .out(wire_253));
  TC_IndexerBit # (.UUID(64'd3061326707059992105 ^ UUID), .INDEX(64'd5)) IndexerBit_306 (.in({{56{1'b0}}, wire_71 }), .out(wire_211));
  TC_Decoder3 # (.UUID(64'd2662776985470781262 ^ UUID)) Decoder3_307 (.dis(wire_292), .sel0(wire_253), .sel1(wire_325), .sel2(wire_211), .out0(wire_78), .out1(wire_352), .out2(wire_124), .out3(wire_109), .out4(wire_177), .out5(wire_297), .out6(), .out7());
  TC_IndexerBit # (.UUID(64'd2678787801262638114 ^ UUID), .INDEX(64'd4)) IndexerBit_308 (.in({{56{1'b0}}, wire_71 }), .out(wire_325));
  TC_Maker8 # (.UUID(64'd3787849024130992586 ^ UUID)) Maker8_309 (.in0(wire_27), .in1(wire_64), .in2(wire_306), .in3(wire_188), .in4(wire_296), .in5(wire_270), .in6(wire_308), .in7(wire_151), .out(wire_313));
  TC_Maker8 # (.UUID(64'd2623625314989675875 ^ UUID)) Maker8_310 (.in0(wire_332), .in1(wire_294), .in2(wire_303), .in3(wire_320), .in4(wire_324), .in5(wire_368), .in6(wire_376), .in7(wire_322), .out(wire_198));
  TC_Maker8 # (.UUID(64'd3386126329111862344 ^ UUID)) Maker8_311 (.in0(wire_240), .in1(wire_104), .in2(wire_360), .in3(wire_102), .in4(wire_231), .in5(wire_384), .in6(wire_365), .in7(wire_184), .out(wire_221));
  TC_Decoder3 # (.UUID(64'd287751819982062857 ^ UUID)) Decoder3_312 (.dis(wire_119[0:0]), .sel0(wire_155[0:0]), .sel1(wire_81[0:0]), .sel2(wire_108[0:0]), .out0(wire_240), .out1(wire_104), .out2(wire_360), .out3(wire_102), .out4(wire_231), .out5(wire_384), .out6(wire_365), .out7(wire_184));
  TC_Decoder3 # (.UUID(64'd798995494482774220 ^ UUID)) Decoder3_313 (.dis(wire_354[0:0]), .sel0(wire_155[0:0]), .sel1(wire_81[0:0]), .sel2(wire_108[0:0]), .out0(wire_332), .out1(wire_294), .out2(wire_303), .out3(wire_320), .out4(wire_324), .out5(wire_368), .out6(wire_376), .out7(wire_322));
  TC_Decoder3 # (.UUID(64'd2575998536381794021 ^ UUID)) Decoder3_314 (.dis(wire_402[0:0]), .sel0(wire_155[0:0]), .sel1(wire_81[0:0]), .sel2(wire_108[0:0]), .out0(wire_27), .out1(wire_64), .out2(wire_306), .out3(wire_188), .out4(wire_296), .out5(wire_270), .out6(wire_308), .out7(wire_151));
  TC_Maker64 # (.UUID(64'd2118416430580755710 ^ UUID)) Maker64_315 (.in0({{7{1'b0}}, wire_23 }), .in1({{7{1'b0}}, wire_138 }), .in2({{7{1'b0}}, wire_30 }), .in3({{7{1'b0}}, wire_247 }), .in4({{7{1'b0}}, wire_128 }), .in5({{7{1'b0}}, wire_142 }), .in6(8'd0), .in7(8'd0), .out(wire_17));
  TC_IndexerByte # (.UUID(64'd4204561175501303620 ^ UUID), .INDEX(64'd0)) IndexerByte_316 (.in(wire_17), .out(wire_155));
  TC_IndexerByte # (.UUID(64'd1496946436106024662 ^ UUID), .INDEX(64'd1)) IndexerByte_317 (.in(wire_17), .out(wire_81));
  TC_IndexerByte # (.UUID(64'd2871709126300377013 ^ UUID), .INDEX(64'd2)) IndexerByte_318 (.in(wire_17), .out(wire_108));
  TC_IndexerByte # (.UUID(64'd3715263176504705704 ^ UUID), .INDEX(64'd3)) IndexerByte_319 (.in(wire_17), .out(wire_119));
  TC_Not # (.UUID(64'd2012876504612309001 ^ UUID), .BIT_WIDTH(64'd1)) Not_320 (.in(wire_297), .out(wire_142));
  TC_Not # (.UUID(64'd2535620781485868088 ^ UUID), .BIT_WIDTH(64'd1)) Not_321 (.in(wire_177), .out(wire_128));
  TC_Not # (.UUID(64'd4486387007616451464 ^ UUID), .BIT_WIDTH(64'd1)) Not_322 (.in(wire_109), .out(wire_247));
  TC_Not # (.UUID(64'd2498440524644937755 ^ UUID), .BIT_WIDTH(64'd1)) Not_323 (.in(wire_124), .out(wire_279));
  TC_Not # (.UUID(64'd336274444425496480 ^ UUID), .BIT_WIDTH(64'd1)) Not_324 (.in(wire_352), .out(wire_374));
  TC_IndexerBit # (.UUID(64'd1121085966967498408 ^ UUID), .INDEX(64'd2)) IndexerBit_325 (.in({{56{1'b0}}, wire_71 }), .out(wire_30));
  TC_IndexerBit # (.UUID(64'd4071184576641035735 ^ UUID), .INDEX(64'd1)) IndexerBit_326 (.in({{56{1'b0}}, wire_71 }), .out(wire_138));
  TC_IndexerBit # (.UUID(64'd1666500121691486869 ^ UUID), .INDEX(64'd0)) IndexerBit_327 (.in({{56{1'b0}}, wire_71 }), .out(wire_23));
  TC_Not # (.UUID(64'd259775706542815838 ^ UUID), .BIT_WIDTH(64'd1)) Not_328 (.in(wire_42), .out(wire_292));
  TC_Maker64 # (.UUID(64'd611788617181826292 ^ UUID)) Maker64_329 (.in0(8'd0), .in1(wire_256), .in2(wire_304), .in3(wire_131), .in4(wire_221), .in5(wire_198), .in6(wire_313), .in7(8'd0), .out(wire_63));
  TC_Switch # (.UUID(64'd552336782343327323 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_330 (.en(wire_42), .in(wire_1[15:0]), .out(wire_318));
  TC_Splitter16 # (.UUID(64'd2056784098263663101 ^ UUID)) Splitter16_331 (.in(wire_318), .out0(wire_193), .out1(wire_52));
  TC_And # (.UUID(64'd4280897558495300328 ^ UUID), .BIT_WIDTH(64'd8)) And8_332 (.in0(wire_52), .in1(wire_175), .out(wire_68));
  TC_Constant # (.UUID(64'd2179588892679277563 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hFC)) Constant8_333 (.out(wire_175));
  TC_Maker16 # (.UUID(64'd4094676674732942649 ^ UUID)) Maker16_334 (.in0(wire_193), .in1(wire_265), .out(wire_202));
  TC_And # (.UUID(64'd553791687166410429 ^ UUID), .BIT_WIDTH(64'd8)) And8_335 (.in0(wire_193), .in1(wire_148), .out(wire_176));
  TC_Constant # (.UUID(64'd2493964338307637551 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1F)) Constant8_336 (.out(wire_148));
  TC_Shr # (.UUID(64'd615409739448528046 ^ UUID), .BIT_WIDTH(64'd16)) Shr16_337 (.in(wire_202), .shift(wire_404), .out(wire_349));
  TC_Mul # (.UUID(64'd2101900763352689865 ^ UUID), .BIT_WIDTH(64'd8)) DivMod8_338 (.in0(wire_349[7:0]), .in1(wire_309), .out0(wire_271), .out1(wire_210));
  TC_And # (.UUID(64'd1530495578126298051 ^ UUID), .BIT_WIDTH(64'd8)) And8_339 (.in0(wire_160), .in1(wire_176), .out(wire_16));
  TC_Shr # (.UUID(64'd4019376895550813305 ^ UUID), .BIT_WIDTH(64'd8)) Shr8_340 (.in(wire_176), .shift(wire_205), .out(wire_249));
  TC_Mul # (.UUID(64'd2508741242317517872 ^ UUID), .BIT_WIDTH(64'd8)) Mul8_341 (.in0(wire_359), .in1(wire_210), .out0(wire_58), .out1());
  TC_Constant # (.UUID(64'd2386342230809029268 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h5)) Constant8_342 (.out(wire_404));
  TC_Add # (.UUID(64'd1080761739701450832 ^ UUID), .BIT_WIDTH(64'd8)) Add8_343 (.in0(wire_58), .in1(wire_16), .ci(1'd0), .out(wire_71), .co());
  TC_Constant # (.UUID(64'd102880999750610880 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h8)) Constant8_344 (.out(wire_359));
  TC_Constant # (.UUID(64'd268383145457663394 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6)) Constant8_345 (.out(wire_309));
  TC_And # (.UUID(64'd3182749074842184933 ^ UUID), .BIT_WIDTH(64'd8)) And8_346 (.in0(wire_52), .in1(wire_375), .out(wire_265));
  TC_Constant # (.UUID(64'd529183091884845671 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7)) Constant8_347 (.out(wire_160));
  TC_Maker16 # (.UUID(64'd3705568547552444440 ^ UUID)) Maker16_348 (.in0(wire_271), .in1(wire_249), .out(wire_39));
  TC_Constant # (.UUID(64'd733594082608262947 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h3)) Constant8_349 (.out(wire_205));
  TC_Constant # (.UUID(64'd755935072730837764 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h3)) Constant8_350 (.out(wire_375));
  TC_IndexerByte # (.UUID(64'd1266734280984969515 ^ UUID), .INDEX(64'd5)) IndexerByte_351 (.in(wire_17), .out(wire_402));
  TC_IndexerByte # (.UUID(64'd3148190672076504148 ^ UUID), .INDEX(64'd4)) IndexerByte_352 (.in(wire_17), .out(wire_354));
  TC_Not # (.UUID(64'd71963519918302721 ^ UUID), .BIT_WIDTH(64'd1)) Not_353 (.in(wire_78), .out(wire_201));
  TC_Equal # (.UUID(64'd2806767944650985817 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_354 (.in0(wire_370), .in1(wire_159), .out(wire_42));
  TC_Constant # (.UUID(64'd3863763634612194638 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hE0)) Constant8_355 (.out(wire_159));
  TC_Splitter16 # (.UUID(64'd1245764572034183129 ^ UUID)) Splitter16_356 (.in(wire_46), .out0(), .out1(wire_370));

  wire [0:0] wire_0;
  wire [63:0] wire_1;
  wire [63:0] wire_1_0;
  wire [63:0] wire_1_1;
  wire [63:0] wire_1_2;
  wire [63:0] wire_1_3;
  wire [63:0] wire_1_4;
  wire [63:0] wire_1_5;
  wire [63:0] wire_1_6;
  wire [63:0] wire_1_7;
  wire [63:0] wire_1_8;
  wire [63:0] wire_1_9;
  wire [63:0] wire_1_10;
  wire [63:0] wire_1_11;
  wire [63:0] wire_1_12;
  wire [63:0] wire_1_13;
  wire [63:0] wire_1_14;
  wire [63:0] wire_1_15;
  wire [63:0] wire_1_16;
  wire [63:0] wire_1_17;
  wire [63:0] wire_1_18;
  wire [63:0] wire_1_19;
  wire [63:0] wire_1_20;
  assign wire_1 = wire_1_0|wire_1_1|wire_1_2|wire_1_3|wire_1_4|wire_1_5|wire_1_6|wire_1_7|wire_1_8|wire_1_9|wire_1_10|wire_1_11|wire_1_12|wire_1_13|wire_1_14|wire_1_15|wire_1_16|wire_1_17|wire_1_18|wire_1_19|wire_1_20;
  wire [0:0] wire_2;
  wire [15:0] wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  wire [7:0] wire_6;
  wire [0:0] wire_7;
  wire [15:0] wire_8;
  wire [31:0] wire_9;
  wire [63:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [15:0] wire_15;
  wire [7:0] wire_16;
  wire [63:0] wire_17;
  wire [0:0] wire_18;
  wire [63:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [31:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [15:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [7:0] wire_34;
  wire [15:0] wire_35;
  wire [15:0] wire_35_0;
  wire [15:0] wire_35_1;
  assign wire_35 = wire_35_0|wire_35_1;
  wire [0:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [15:0] wire_39;
  wire [0:0] wire_40;
  wire [7:0] wire_41;
  wire [0:0] wire_42;
  wire [15:0] wire_43;
  wire [0:0] wire_44;
  wire [15:0] wire_45;
  wire [15:0] wire_46;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  wire [0:0] wire_49;
  wire [63:0] wire_50;
  wire [0:0] wire_51;
  wire [7:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  wire [0:0] wire_54_0;
  wire [0:0] wire_54_1;
  wire [0:0] wire_54_2;
  wire [0:0] wire_54_3;
  wire [0:0] wire_54_4;
  wire [0:0] wire_54_5;
  wire [0:0] wire_54_6;
  wire [0:0] wire_54_7;
  wire [0:0] wire_54_8;
  wire [0:0] wire_54_9;
  assign wire_54 = wire_54_0|wire_54_1|wire_54_2|wire_54_3|wire_54_4|wire_54_5|wire_54_6|wire_54_7|wire_54_8|wire_54_9;
  wire [0:0] wire_55;
  wire [31:0] wire_56;
  wire [7:0] wire_57;
  wire [7:0] wire_58;
  wire [0:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [15:0] wire_62;
  wire [63:0] wire_63;
  wire [0:0] wire_64;
  wire [0:0] wire_65;
  wire [15:0] wire_66;
  wire [0:0] wire_67;
  wire [7:0] wire_68;
  wire [0:0] wire_69;
  wire [0:0] wire_70;
  wire [7:0] wire_71;
  wire [0:0] wire_72;
  wire [0:0] wire_73;
  wire [15:0] wire_74;
  wire [0:0] wire_75;
  wire [0:0] wire_76;
  wire [0:0] wire_77;
  wire [0:0] wire_78;
  wire [0:0] wire_79;
  wire [0:0] wire_80;
  wire [7:0] wire_81;
  wire [0:0] wire_82;
  wire [63:0] wire_83;
  wire [15:0] wire_84;
  wire [15:0] wire_85;
  wire [15:0] wire_86;
  wire [0:0] wire_87;
  wire [0:0] wire_88;
  wire [7:0] wire_89;
  wire [0:0] wire_90;
  wire [0:0] wire_91;
  wire [0:0] wire_92;
  assign arch_output_enable = wire_92;
  wire [0:0] wire_93;
  wire [0:0] wire_94;
  wire [0:0] wire_95;
  wire [7:0] wire_96;
  wire [15:0] wire_97;
  wire [15:0] wire_97_0;
  wire [15:0] wire_97_1;
  assign wire_97 = wire_97_0|wire_97_1;
  wire [15:0] wire_98;
  wire [15:0] wire_98_0;
  wire [15:0] wire_98_1;
  assign wire_98 = wire_98_0|wire_98_1;
  wire [0:0] wire_99;
  wire [7:0] wire_100;
  wire [31:0] wire_101;
  wire [0:0] wire_102;
  wire [0:0] wire_103;
  wire [0:0] wire_104;
  wire [0:0] wire_105;
  wire [7:0] wire_106;
  wire [0:0] wire_107;
  wire [7:0] wire_108;
  wire [0:0] wire_109;
  wire [7:0] wire_110;
  wire [0:0] wire_111;
  wire [0:0] wire_112;
  wire [0:0] wire_113;
  wire [0:0] wire_114;
  wire [0:0] wire_115;
  wire [7:0] wire_116;
  wire [15:0] wire_117;
  wire [0:0] wire_118;
  wire [7:0] wire_119;
  wire [0:0] wire_120;
  wire [0:0] wire_121;
  wire [7:0] wire_122;
  wire [7:0] wire_123;
  wire [0:0] wire_124;
  wire [15:0] wire_125;
  wire [63:0] wire_126;
  wire [15:0] wire_127;
  wire [15:0] wire_127_0;
  wire [15:0] wire_127_1;
  assign wire_127 = wire_127_0|wire_127_1;
  wire [0:0] wire_128;
  wire [7:0] wire_129;
  wire [0:0] wire_130;
  wire [7:0] wire_131;
  wire [15:0] wire_132;
  wire [0:0] wire_133;
  wire [7:0] wire_134;
  wire [0:0] wire_135;
  wire [15:0] wire_136;
  wire [15:0] wire_136_0;
  wire [15:0] wire_136_1;
  wire [15:0] wire_136_2;
  assign wire_136 = wire_136_0|wire_136_1|wire_136_2;
  wire [7:0] wire_137;
  wire [0:0] wire_138;
  wire [31:0] wire_139;
  wire [0:0] wire_140;
  wire [7:0] wire_141;
  wire [0:0] wire_142;
  wire [63:0] wire_143;
  wire [15:0] wire_144;
  wire [0:0] wire_145;
  wire [0:0] wire_146;
  wire [15:0] wire_147;
  wire [7:0] wire_148;
  wire [15:0] wire_149;
  wire [7:0] wire_150;
  wire [0:0] wire_151;
  wire [15:0] wire_152;
  wire [63:0] wire_153;
  wire [0:0] wire_154;
  wire [7:0] wire_155;
  wire [0:0] wire_156;
  wire [0:0] wire_157;
  wire [7:0] wire_158;
  wire [7:0] wire_159;
  wire [7:0] wire_160;
  wire [15:0] wire_161;
  wire [0:0] wire_162;
  wire [0:0] wire_163;
  wire [0:0] wire_164;
  wire [63:0] wire_165;
  wire [0:0] wire_166;
  wire [15:0] wire_167;
  wire [7:0] wire_168;
  wire [63:0] wire_169;
  wire [0:0] wire_170;
  wire [0:0] wire_171;
  wire [15:0] wire_172;
  wire [7:0] wire_173;
  wire [0:0] wire_174;
  wire [7:0] wire_175;
  wire [7:0] wire_176;
  wire [0:0] wire_177;
  wire [31:0] wire_178;
  wire [15:0] wire_179;
  wire [0:0] wire_180;
  wire [15:0] wire_181;
  wire [0:0] wire_182;
  wire [0:0] wire_183;
  wire [0:0] wire_184;
  wire [15:0] wire_185;
  wire [0:0] wire_186;
  wire [63:0] wire_187;
  wire [0:0] wire_188;
  wire [15:0] wire_189;
  wire [15:0] wire_190;
  wire [63:0] wire_191;
  wire [0:0] wire_192;
  wire [7:0] wire_193;
  wire [0:0] wire_194;
  wire [0:0] wire_195;
  wire [0:0] wire_196;
  wire [0:0] wire_197;
  wire [7:0] wire_198;
  wire [0:0] wire_199;
  wire [0:0] wire_200;
  wire [0:0] wire_201;
  wire [15:0] wire_202;
  wire [15:0] wire_203;
  wire [15:0] wire_204;
  wire [7:0] wire_205;
  wire [0:0] wire_206;
  wire [0:0] wire_207;
  wire [7:0] wire_208;
  wire [0:0] wire_209;
  wire [7:0] wire_210;
  wire [0:0] wire_211;
  wire [0:0] wire_212;
  wire [0:0] wire_213;
  wire [0:0] wire_214;
  wire [0:0] wire_214_0;
  wire [0:0] wire_214_1;
  wire [0:0] wire_214_2;
  assign wire_214 = wire_214_0|wire_214_1|wire_214_2;
  wire [0:0] wire_215;
  wire [0:0] wire_216;
  wire [63:0] wire_217;
  wire [63:0] wire_218;
  wire [31:0] wire_219;
  wire [0:0] wire_220;
  wire [7:0] wire_221;
  wire [0:0] wire_222;
  wire [0:0] wire_223;
  wire [0:0] wire_224;
  wire [7:0] wire_225;
  wire [0:0] wire_226;
  wire [0:0] wire_227;
  wire [7:0] wire_228;
  wire [0:0] wire_229;
  wire [0:0] wire_230;
  wire [0:0] wire_231;
  wire [0:0] wire_232;
  wire [7:0] wire_233;
  wire [0:0] wire_234;
  wire [15:0] wire_235;
  wire [7:0] wire_236;
  wire [0:0] wire_237;
  wire [0:0] wire_238;
  wire [15:0] wire_239;
  wire [0:0] wire_240;
  wire [7:0] wire_241;
  wire [15:0] wire_242;
  wire [0:0] wire_243;
  wire [31:0] wire_244;
  wire [0:0] wire_245;
  wire [0:0] wire_246;
  wire [0:0] wire_247;
  wire [63:0] wire_248;
  wire [7:0] wire_249;
  wire [63:0] wire_250;
  wire [0:0] wire_251;
  wire [0:0] wire_252;
  wire [0:0] wire_253;
  wire [0:0] wire_254;
  wire [0:0] wire_255;
  wire [7:0] wire_256;
  wire [0:0] wire_257;
  wire [0:0] wire_258;
  wire [0:0] wire_259;
  wire [0:0] wire_260;
  wire [0:0] wire_261;
  wire [0:0] wire_262;
  wire [15:0] wire_263;
  wire [0:0] wire_264;
  wire [7:0] wire_265;
  wire [0:0] wire_266;
  wire [0:0] wire_267;
  wire [0:0] wire_268;
  wire [15:0] wire_269;
  wire [0:0] wire_270;
  wire [7:0] wire_271;
  wire [0:0] wire_272;
  wire [0:0] wire_273;
  wire [7:0] wire_274;
  wire [7:0] wire_275;
  wire [0:0] wire_276;
  wire [0:0] wire_277;
  wire [7:0] wire_278;
  wire [0:0] wire_279;
  wire [15:0] wire_280;
  wire [0:0] wire_281;
  wire [15:0] wire_282;
  wire [15:0] wire_283;
  wire [0:0] wire_284;
  wire [15:0] wire_285;
  wire [15:0] wire_286;
  wire [0:0] wire_287;
  wire [0:0] wire_288;
  wire [0:0] wire_289;
  wire [63:0] wire_290;
  wire [7:0] wire_291;
  wire [0:0] wire_292;
  wire [7:0] wire_293;
  wire [0:0] wire_294;
  wire [0:0] wire_295;
  wire [0:0] wire_296;
  wire [0:0] wire_297;
  wire [0:0] wire_298;
  wire [0:0] wire_299;
  wire [0:0] wire_300;
  wire [0:0] wire_301;
  wire [0:0] wire_302;
  wire [0:0] wire_303;
  wire [7:0] wire_304;
  wire [15:0] wire_305;
  wire [0:0] wire_306;
  wire [15:0] wire_307;
  wire [0:0] wire_308;
  wire [7:0] wire_309;
  wire [0:0] wire_310;
  wire [0:0] wire_311;
  wire [15:0] wire_312;
  wire [7:0] wire_313;
  wire [0:0] wire_314;
  wire [0:0] wire_315;
  wire [0:0] wire_316;
  wire [0:0] wire_317;
  wire [15:0] wire_318;
  wire [0:0] wire_319;
  wire [0:0] wire_320;
  wire [0:0] wire_321;
  wire [0:0] wire_322;
  wire [7:0] wire_323;
  wire [0:0] wire_324;
  wire [0:0] wire_325;
  wire [0:0] wire_326;
  wire [0:0] wire_327;
  wire [7:0] wire_328;
  wire [0:0] wire_329;
  wire [0:0] wire_330;
  wire [0:0] wire_331;
  wire [0:0] wire_332;
  wire [0:0] wire_333;
  wire [0:0] wire_334;
  wire [0:0] wire_335;
  assign arch_input_enable = wire_335;
  wire [15:0] wire_336;
  wire [0:0] wire_337;
  wire [0:0] wire_338;
  wire [0:0] wire_339;
  wire [7:0] wire_340;
  wire [15:0] wire_341;
  wire [0:0] wire_342;
  wire [0:0] wire_343;
  wire [0:0] wire_344;
  wire [0:0] wire_345;
  wire [7:0] wire_346;
  wire [7:0] wire_347;
  wire [7:0] wire_348;
  wire [15:0] wire_349;
  wire [0:0] wire_350;
  wire [0:0] wire_351;
  wire [0:0] wire_352;
  wire [0:0] wire_353;
  wire [7:0] wire_354;
  wire [0:0] wire_355;
  wire [0:0] wire_356;
  wire [0:0] wire_357;
  wire [0:0] wire_358;
  wire [7:0] wire_359;
  wire [0:0] wire_360;
  wire [15:0] wire_361;
  wire [0:0] wire_362;
  wire [0:0] wire_363;
  wire [0:0] wire_364;
  assign wire_364 = 0;
  wire [0:0] wire_365;
  wire [0:0] wire_366;
  wire [0:0] wire_367;
  wire [0:0] wire_368;
  wire [15:0] wire_369;
  wire [7:0] wire_370;
  wire [0:0] wire_371;
  wire [0:0] wire_372;
  wire [7:0] wire_373;
  wire [0:0] wire_374;
  wire [7:0] wire_375;
  wire [0:0] wire_376;
  wire [0:0] wire_377;
  wire [0:0] wire_378;
  wire [63:0] wire_379;
  wire [0:0] wire_380;
  wire [63:0] wire_381;
  wire [0:0] wire_382;
  wire [15:0] wire_383;
  wire [0:0] wire_384;
  wire [0:0] wire_385;
  wire [63:0] wire_386;
  wire [15:0] wire_387;
  wire [15:0] wire_388;
  wire [0:0] wire_389;
  wire [7:0] wire_390;
  wire [0:0] wire_391;
  wire [0:0] wire_392;
  wire [0:0] wire_393;
  wire [0:0] wire_394;
  wire [0:0] wire_395;
  wire [0:0] wire_396;
  wire [0:0] wire_397;
  wire [7:0] wire_398;
  wire [7:0] wire_399;
  wire [15:0] wire_400;
  wire [15:0] wire_401;
  wire [7:0] wire_402;
  wire [15:0] wire_403;
  wire [7:0] wire_404;
  wire [0:0] wire_405;
  wire [0:0] wire_406;
  wire [15:0] wire_407;
  wire [0:0] wire_408;
  wire [0:0] wire_409;

endmodule
